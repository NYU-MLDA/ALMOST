//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n202_), .A3(KEYINPUT21), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT85), .ZN(new_n213_));
  INV_X1    g012(.A(G155gat), .ZN(new_n214_));
  INV_X1    g013(.A(G162gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(KEYINPUT86), .B2(KEYINPUT3), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT87), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n219_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n221_), .A2(KEYINPUT86), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT84), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n224_), .A2(new_n227_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n218_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n217_), .A2(KEYINPUT1), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n216_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n213_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n225_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n211_), .B1(new_n243_), .B2(KEYINPUT29), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G228gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(KEYINPUT88), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(KEYINPUT88), .ZN(new_n249_));
  XOR2_X1   g048(.A(G78gat), .B(G106gat), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n243_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT28), .B1(new_n243_), .B2(KEYINPUT29), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G22gat), .B(G50gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n249_), .A2(new_n251_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n251_), .B1(new_n249_), .B2(new_n259_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n248_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n249_), .A2(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n250_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n247_), .A3(new_n260_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(G85gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT0), .B(G57gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n218_), .A2(new_n235_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G127gat), .B(G134gat), .Z(new_n274_));
  XOR2_X1   g073(.A(G113gat), .B(G120gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n273_), .A2(KEYINPUT4), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n236_), .A2(new_n281_), .A3(new_n242_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT93), .A3(new_n276_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n276_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n243_), .B2(KEYINPUT93), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n273_), .B2(new_n281_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n283_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT4), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT95), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(KEYINPUT95), .A3(KEYINPUT4), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n280_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n278_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n272_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n282_), .A2(KEYINPUT93), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n276_), .B1(new_n273_), .B2(new_n286_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI211_X1 g099(.A(new_n290_), .B(new_n297_), .C1(new_n300_), .C2(new_n283_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT95), .B1(new_n288_), .B2(KEYINPUT4), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n279_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(new_n294_), .A3(new_n271_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(KEYINPUT98), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT98), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n306_), .B(new_n272_), .C1(new_n293_), .C2(new_n295_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT27), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT91), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT22), .B(G169gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT90), .ZN(new_n320_));
  INV_X1    g119(.A(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(KEYINPUT91), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n317_), .A2(new_n318_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G190gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT89), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT25), .B(G183gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n329_), .A2(KEYINPUT24), .A3(new_n318_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(KEYINPUT24), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n330_), .A2(new_n314_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n211_), .B1(new_n324_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n327_), .A2(new_n325_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G169gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT20), .B1(new_n340_), .B2(new_n210_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n311_), .B1(new_n334_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n324_), .A2(new_n211_), .A3(new_n333_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n311_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n210_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n343_), .A2(KEYINPUT20), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G8gat), .B(G36gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n309_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n352_), .B(KEYINPUT99), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n343_), .A2(KEYINPUT20), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT97), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT97), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n343_), .A2(new_n360_), .A3(KEYINPUT20), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n345_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n311_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n334_), .A2(new_n341_), .A3(new_n311_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n357_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT100), .B1(new_n347_), .B2(new_n353_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT100), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n342_), .A2(new_n346_), .A3(new_n368_), .A4(new_n352_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(KEYINPUT27), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n356_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G71gat), .B(G99gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G43gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n340_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(new_n284_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(G15gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT30), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT31), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n376_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n267_), .A2(new_n308_), .A3(new_n372_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n304_), .A2(KEYINPUT96), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT33), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n304_), .A2(KEYINPUT96), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n354_), .A2(new_n355_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n278_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n277_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n271_), .B1(new_n288_), .B2(new_n390_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n389_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n386_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n364_), .B1(new_n362_), .B2(new_n311_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n397_));
  MUX2_X1   g196(.A(new_n396_), .B(new_n347_), .S(new_n397_), .Z(new_n398_));
  NAND3_X1  g197(.A1(new_n305_), .A2(new_n307_), .A3(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n395_), .A2(new_n267_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n371_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n382_), .B1(new_n401_), .B2(new_n267_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n384_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT73), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G85gat), .A2(G92gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(G85gat), .A2(G92gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(KEYINPUT9), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT64), .B(G85gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT65), .B(G92gat), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n407_), .B1(new_n410_), .B2(KEYINPUT9), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G99gat), .A2(G106gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT6), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(G99gat), .A3(G106gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G106gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT10), .B(G99gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n411_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G71gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT69), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G71gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(G78gat), .ZN(new_n427_));
  INV_X1    g226(.A(G78gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G64gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G57gat), .ZN(new_n431_));
  INV_X1    g230(.A(G57gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G64gat), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n431_), .A2(new_n433_), .A3(KEYINPUT11), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT11), .B1(new_n431_), .B2(new_n433_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n427_), .B(new_n429_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n433_), .A3(KEYINPUT11), .ZN(new_n437_));
  INV_X1    g236(.A(new_n429_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n428_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT8), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n413_), .A2(new_n415_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT67), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n450_));
  INV_X1    g249(.A(G99gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n417_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(KEYINPUT68), .A3(new_n446_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n413_), .A2(new_n415_), .A3(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n444_), .A2(new_n449_), .A3(new_n453_), .A4(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n406_), .A2(new_n405_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n442_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n442_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n452_), .A2(new_n446_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT66), .B1(new_n416_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n447_), .A2(new_n448_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n443_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n459_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n421_), .B(new_n441_), .C1(new_n458_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT72), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n421_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT70), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n459_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n416_), .A2(new_n460_), .A3(KEYINPUT66), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n463_), .B1(new_n462_), .B2(new_n443_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n457_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n452_), .A2(KEYINPUT68), .A3(new_n446_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT68), .B1(new_n452_), .B2(new_n446_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n413_), .A2(new_n415_), .A3(new_n454_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n454_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n479_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n478_), .B(KEYINPUT70), .C1(new_n486_), .C2(new_n442_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n472_), .B1(new_n474_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n441_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT12), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n478_), .B1(new_n486_), .B2(new_n442_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n441_), .B1(new_n491_), .B2(new_n421_), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI22_X1  g293(.A1(new_n488_), .A2(new_n490_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n404_), .B1(new_n471_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n466_), .A2(new_n468_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT72), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n490_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n474_), .A2(new_n487_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n472_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n458_), .A2(new_n465_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n472_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n493_), .B1(new_n505_), .B2(new_n441_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n500_), .A2(new_n503_), .A3(KEYINPUT73), .A4(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n468_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n466_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n492_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n496_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G120gat), .B(G148gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT5), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G176gat), .B(G204gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n496_), .A2(new_n507_), .A3(new_n510_), .A4(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(KEYINPUT74), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT74), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n511_), .A2(new_n520_), .A3(new_n515_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n519_), .A2(KEYINPUT13), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT13), .B1(new_n519_), .B2(new_n521_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G36gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(G29gat), .ZN(new_n528_));
  INV_X1    g327(.A(G29gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G36gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n530_), .A3(KEYINPUT77), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT77), .B1(new_n528_), .B2(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n526_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n530_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT77), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(new_n531_), .A3(new_n525_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n538_), .A3(KEYINPUT15), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543_));
  INV_X1    g342(.A(G1gat), .ZN(new_n544_));
  INV_X1    g343(.A(G8gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G8gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT83), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n532_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n525_), .B1(new_n537_), .B2(new_n531_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n547_), .B(new_n548_), .Z(new_n555_));
  NAND3_X1  g354(.A1(new_n534_), .A2(new_n538_), .A3(KEYINPUT83), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n534_), .A2(KEYINPUT83), .A3(new_n538_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT83), .B1(new_n534_), .B2(new_n538_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n549_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n555_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n559_), .B1(new_n564_), .B2(new_n558_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n565_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n524_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n403_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT35), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n505_), .B2(new_n539_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n541_), .A2(new_n542_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n488_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(KEYINPUT35), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT76), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n578_), .B(new_n582_), .C1(new_n488_), .C2(new_n579_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT36), .Z(new_n590_));
  AND2_X1   g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT78), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n584_), .A2(new_n585_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n591_), .A2(new_n596_), .A3(KEYINPUT37), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n586_), .A2(new_n590_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT80), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT79), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n584_), .A2(KEYINPUT79), .A3(new_n585_), .A4(new_n594_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n586_), .A2(KEYINPUT80), .A3(new_n590_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .A4(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n597_), .B1(new_n605_), .B2(KEYINPUT37), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n549_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n441_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT81), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n610_), .A2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n616_), .B2(new_n614_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n609_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n606_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT82), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n573_), .A2(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n625_), .A2(G1gat), .A3(new_n308_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n598_), .A2(KEYINPUT101), .A3(new_n595_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT101), .B1(new_n598_), .B2(new_n595_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n308_), .A2(new_n372_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n263_), .A2(new_n266_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n395_), .A2(new_n267_), .A3(new_n399_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n382_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n630_), .B1(new_n635_), .B2(new_n384_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n621_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n572_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n308_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n544_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT38), .B1(new_n626_), .B2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(KEYINPUT38), .B2(new_n626_), .ZN(G1324gat));
  INV_X1    g441(.A(new_n625_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n545_), .A3(new_n371_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT102), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n545_), .B1(new_n638_), .B2(new_n371_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(KEYINPUT40), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  AOI21_X1  g452(.A(new_n378_), .B1(new_n638_), .B2(new_n383_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n643_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(G22gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n638_), .B2(new_n632_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n643_), .A2(new_n658_), .A3(new_n632_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  NOR2_X1   g462(.A1(new_n629_), .A2(new_n637_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n573_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n639_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n403_), .A2(new_n606_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT43), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n403_), .A2(new_n669_), .A3(new_n606_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n572_), .A2(new_n621_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n671_), .A2(KEYINPUT44), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT44), .B1(new_n671_), .B2(new_n673_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n308_), .A2(new_n529_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n666_), .B1(new_n676_), .B2(new_n677_), .ZN(G1328gat));
  NAND3_X1  g477(.A1(new_n665_), .A2(new_n527_), .A3(new_n371_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT45), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n674_), .A2(new_n675_), .A3(new_n372_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n527_), .B2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI221_X1 g483(.A(new_n680_), .B1(KEYINPUT104), .B2(KEYINPUT46), .C1(new_n527_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1329gat));
  AOI21_X1  g485(.A(G43gat), .B1(new_n665_), .B2(new_n383_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n383_), .A2(G43gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n676_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1330gat));
  INV_X1    g490(.A(G50gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n665_), .A2(new_n692_), .A3(new_n632_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n676_), .A2(new_n694_), .A3(new_n632_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n676_), .B2(new_n632_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1331gat));
  NOR3_X1   g497(.A1(new_n522_), .A2(new_n523_), .A3(new_n570_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n403_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n624_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n432_), .A3(new_n639_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n699_), .A2(new_n637_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n636_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n308_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(G1332gat));
  OAI21_X1  g505(.A(G64gat), .B1(new_n704_), .B2(new_n372_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT48), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n701_), .A2(new_n430_), .A3(new_n371_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  NOR2_X1   g509(.A1(new_n382_), .A2(G71gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT107), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n701_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n704_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n383_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT106), .B(KEYINPUT49), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(G71gat), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n715_), .B2(G71gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT108), .Z(G1334gat));
  NAND3_X1  g519(.A1(new_n701_), .A2(new_n428_), .A3(new_n632_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G78gat), .B1(new_n704_), .B2(new_n267_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT50), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT50), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT109), .ZN(G1335gat));
  NAND2_X1  g525(.A1(new_n605_), .A2(KEYINPUT37), .ZN(new_n727_));
  INV_X1    g526(.A(new_n597_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT43), .B(new_n729_), .C1(new_n635_), .C2(new_n384_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n669_), .B1(new_n403_), .B2(new_n606_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n671_), .A2(KEYINPUT110), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n699_), .A2(new_n621_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n639_), .A2(new_n408_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n700_), .A2(new_n664_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n639_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1336gat));
  AOI21_X1  g540(.A(G92gat), .B1(new_n739_), .B2(new_n371_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT111), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n371_), .A2(new_n409_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n735_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1337gat));
  NOR3_X1   g545(.A1(new_n738_), .A2(new_n418_), .A3(new_n382_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n732_), .A2(new_n733_), .A3(new_n383_), .A4(new_n734_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G99gat), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT51), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT113), .Z(new_n752_));
  XOR2_X1   g551(.A(new_n749_), .B(new_n752_), .Z(G1338gat));
  NAND3_X1  g552(.A1(new_n739_), .A2(new_n417_), .A3(new_n632_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n699_), .A2(new_n632_), .A3(new_n621_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n757_), .B(KEYINPUT114), .C1(new_n730_), .C2(new_n731_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n417_), .B1(new_n755_), .B2(KEYINPUT52), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n756_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n756_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n763_), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n765_), .B(new_n766_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n754_), .B1(new_n764_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n770_), .B(new_n754_), .C1(new_n764_), .C2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  INV_X1    g573(.A(new_n558_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n549_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n557_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT117), .B1(new_n777_), .B2(new_n568_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n558_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n569_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n550_), .A2(new_n557_), .A3(new_n775_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT118), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n565_), .A2(new_n569_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n783_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n518_), .A2(new_n785_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT119), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n518_), .A2(new_n790_), .A3(new_n785_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n496_), .A2(new_n507_), .A3(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT116), .B(new_n508_), .C1(new_n495_), .C2(new_n509_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n500_), .A2(new_n503_), .A3(KEYINPUT55), .A4(new_n506_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n508_), .B1(new_n495_), .B2(new_n509_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .A4(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n515_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n515_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n795_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n729_), .B1(new_n774_), .B2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n795_), .B(KEYINPUT58), .C1(new_n804_), .C2(new_n805_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n518_), .A2(new_n570_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n802_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n496_), .A2(new_n796_), .A3(new_n507_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n515_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n515_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n809_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AND4_X1   g615(.A1(new_n521_), .A2(new_n519_), .A3(new_n785_), .A4(new_n790_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n629_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n807_), .A2(new_n808_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT57), .B(new_n629_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n637_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n729_), .A2(new_n637_), .A3(new_n571_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT54), .B1(new_n823_), .B2(new_n524_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n524_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n622_), .A3(new_n826_), .A4(new_n571_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n773_), .B1(new_n822_), .B2(new_n829_), .ZN(new_n830_));
  NOR4_X1   g629(.A1(new_n308_), .A2(new_n632_), .A3(new_n371_), .A4(new_n382_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n818_), .A2(new_n819_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n806_), .A2(new_n774_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n606_), .A3(new_n808_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n834_), .A3(new_n821_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n621_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(KEYINPUT120), .A3(new_n828_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n830_), .A2(new_n831_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n835_), .A2(new_n842_), .A3(new_n621_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n829_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n831_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n840_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n835_), .A2(new_n842_), .A3(new_n621_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n842_), .B1(new_n835_), .B2(new_n621_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n828_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT122), .A3(new_n845_), .A4(new_n831_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n839_), .A2(new_n847_), .A3(new_n570_), .A4(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G113gat), .ZN(new_n853_));
  OR3_X1    g652(.A1(new_n838_), .A2(G113gat), .A3(new_n571_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1340gat));
  NAND4_X1  g654(.A1(new_n839_), .A2(new_n847_), .A3(new_n524_), .A4(new_n851_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G120gat), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n830_), .A2(new_n837_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n825_), .A2(KEYINPUT60), .ZN(new_n859_));
  MUX2_X1   g658(.A(new_n859_), .B(KEYINPUT60), .S(G120gat), .Z(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n831_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n861_), .ZN(G1341gat));
  NOR2_X1   g661(.A1(new_n621_), .A2(KEYINPUT123), .ZN(new_n863_));
  MUX2_X1   g662(.A(KEYINPUT123), .B(new_n863_), .S(G127gat), .Z(new_n864_));
  NAND4_X1  g663(.A1(new_n839_), .A2(new_n847_), .A3(new_n851_), .A4(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G127gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n838_), .B2(new_n621_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1342gat));
  INV_X1    g667(.A(G134gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n729_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n839_), .A2(new_n847_), .A3(new_n851_), .A4(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n838_), .B2(new_n629_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT124), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n874_), .B(new_n869_), .C1(new_n838_), .C2(new_n629_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n871_), .A2(new_n873_), .A3(new_n875_), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n267_), .A2(new_n383_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n878_), .A2(new_n308_), .A3(new_n371_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n858_), .A2(new_n570_), .A3(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n858_), .A2(new_n524_), .A3(new_n879_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g682(.A1(new_n858_), .A2(new_n637_), .A3(new_n879_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  NAND2_X1  g685(.A1(new_n858_), .A2(new_n879_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G162gat), .B1(new_n887_), .B2(new_n729_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n630_), .A2(new_n215_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(G1347gat));
  NAND3_X1  g689(.A1(new_n308_), .A2(new_n371_), .A3(new_n383_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n632_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n850_), .A2(new_n570_), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n893_), .A2(new_n894_), .A3(G169gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n850_), .A2(new_n892_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(new_n320_), .A3(new_n570_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n893_), .B2(G169gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n895_), .B1(new_n898_), .B2(new_n899_), .ZN(G1348gat));
  AOI21_X1  g699(.A(G176gat), .B1(new_n897_), .B2(new_n524_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n858_), .A2(new_n267_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n825_), .A2(new_n321_), .A3(new_n891_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NOR3_X1   g703(.A1(new_n896_), .A2(new_n327_), .A3(new_n621_), .ZN(new_n905_));
  INV_X1    g704(.A(G183gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n891_), .A2(new_n621_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n858_), .A2(new_n267_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n906_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n896_), .B2(new_n729_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n630_), .A2(new_n326_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n896_), .B2(new_n911_), .ZN(G1351gat));
  NOR3_X1   g711(.A1(new_n878_), .A2(new_n639_), .A3(new_n372_), .ZN(new_n913_));
  OR2_X1    g712(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n914_));
  AND4_X1   g713(.A1(new_n570_), .A2(new_n858_), .A3(new_n913_), .A4(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n858_), .A2(new_n570_), .A3(new_n913_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT125), .B(G197gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1352gat));
  NAND3_X1  g717(.A1(new_n858_), .A2(new_n524_), .A3(new_n913_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n921_));
  INV_X1    g720(.A(G211gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n637_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT126), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n858_), .A2(new_n913_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n922_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1354gat));
  NAND4_X1  g726(.A1(new_n830_), .A2(new_n606_), .A3(new_n837_), .A4(new_n913_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G218gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n629_), .A2(G218gat), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n830_), .A2(new_n837_), .A3(new_n913_), .A4(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT127), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n929_), .A2(new_n934_), .A3(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1355gat));
endmodule


