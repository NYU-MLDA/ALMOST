//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n203_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT25), .B(G183gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT77), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n204_), .B1(G169gat), .B2(G176gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n208_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n211_), .A2(KEYINPUT77), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n205_), .A2(KEYINPUT78), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n205_), .A2(KEYINPUT78), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT22), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(G176gat), .B1(new_n219_), .B2(KEYINPUT79), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(KEYINPUT79), .C2(new_n219_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n203_), .A2(new_n223_), .B1(G169gat), .B2(G176gat), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n215_), .A2(new_n216_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226_));
  OR2_X1    g025(.A1(G127gat), .A2(G134gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G127gat), .A2(G134gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G113gat), .ZN(new_n230_));
  INV_X1    g029(.A(G113gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n231_), .A3(new_n228_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(G120gat), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(G120gat), .B1(new_n230_), .B2(new_n232_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n226_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n232_), .ZN(new_n237_));
  INV_X1    g036(.A(G120gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(KEYINPUT81), .A3(new_n233_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n225_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G99gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT31), .ZN(new_n247_));
  XOR2_X1   g046(.A(G15gat), .B(G43gat), .Z(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  NAND2_X1  g050(.A1(new_n242_), .A2(new_n243_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n245_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n245_), .B2(new_n252_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT90), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G22gat), .B(G50gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT28), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT82), .Z(new_n262_));
  INV_X1    g061(.A(KEYINPUT83), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(G155gat), .B2(G162gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT1), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n270_), .A3(KEYINPUT83), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(KEYINPUT1), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n260_), .B(new_n262_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n261_), .B(KEYINPUT3), .Z(new_n275_));
  XOR2_X1   g074(.A(new_n260_), .B(KEYINPUT2), .Z(new_n276_));
  OAI211_X1 g075(.A(new_n269_), .B(new_n268_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n259_), .B1(new_n278_), .B2(KEYINPUT29), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n274_), .A2(new_n280_), .A3(new_n277_), .A4(new_n258_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n284_));
  XOR2_X1   g083(.A(G211gat), .B(G218gat), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G197gat), .ZN(new_n288_));
  INV_X1    g087(.A(G197gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n288_), .A2(new_n290_), .A3(new_n291_), .A4(KEYINPUT21), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT85), .B1(new_n289_), .B2(G204gat), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n294_), .A2(KEYINPUT21), .B1(new_n288_), .B2(new_n290_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n286_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT86), .B(new_n286_), .C1(new_n293_), .C2(new_n295_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n288_), .A2(new_n290_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n285_), .A2(KEYINPUT21), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT87), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT87), .ZN(new_n304_));
  INV_X1    g103(.A(new_n302_), .ZN(new_n305_));
  AOI211_X1 g104(.A(new_n304_), .B(new_n305_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n283_), .B(new_n284_), .C1(new_n303_), .C2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G78gat), .B(G106gat), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT88), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n294_), .A2(KEYINPUT21), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n301_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n292_), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT86), .B1(new_n314_), .B2(new_n286_), .ZN(new_n315_));
  AOI211_X1 g114(.A(new_n297_), .B(new_n285_), .C1(new_n313_), .C2(new_n292_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n302_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n284_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n283_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n307_), .A2(new_n311_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n311_), .B1(new_n307_), .B2(new_n320_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n282_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT89), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n325_), .B(new_n282_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n307_), .A2(new_n309_), .A3(new_n320_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n309_), .B1(new_n307_), .B2(new_n320_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n279_), .A2(KEYINPUT84), .A3(new_n281_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT84), .B1(new_n279_), .B2(new_n281_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n328_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n256_), .B1(new_n327_), .B2(new_n334_), .ZN(new_n335_));
  AOI211_X1 g134(.A(KEYINPUT90), .B(new_n333_), .C1(new_n324_), .C2(new_n326_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n255_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n307_), .A2(new_n320_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n310_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n307_), .A2(new_n311_), .A3(new_n320_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n325_), .B1(new_n341_), .B2(new_n282_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n326_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n334_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT90), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n327_), .A2(new_n256_), .A3(new_n334_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n255_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT0), .B(G57gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G85gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(G1gat), .B(G29gat), .Z(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n236_), .A2(new_n240_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n234_), .A2(new_n235_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n355_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT4), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT4), .B1(new_n241_), .B2(new_n278_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n241_), .A2(new_n278_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n353_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n352_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n352_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n362_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n358_), .B1(new_n367_), .B2(KEYINPUT4), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n363_), .B(new_n366_), .C1(new_n368_), .C2(new_n353_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n369_), .A3(KEYINPUT93), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT93), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n371_), .B(new_n352_), .C1(new_n360_), .C2(new_n364_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n337_), .A2(new_n348_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n317_), .A2(new_n304_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n300_), .A2(KEYINPUT87), .A3(new_n302_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n225_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT20), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT91), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n224_), .B1(G176gat), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n208_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n317_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n378_), .A2(new_n390_), .A3(KEYINPUT20), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n380_), .A2(new_n382_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n303_), .A2(new_n306_), .ZN(new_n393_));
  OAI221_X1 g192(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n388_), .C1(new_n393_), .C2(new_n225_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n382_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n392_), .A2(new_n402_), .A3(new_n396_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(KEYINPUT27), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n380_), .A2(new_n395_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n394_), .A2(new_n382_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n402_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT95), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT27), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n403_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT95), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n416_), .A3(new_n404_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT96), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n411_), .A2(KEYINPUT95), .B1(new_n403_), .B2(new_n397_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n416_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n407_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n335_), .A2(new_n336_), .A3(new_n255_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n410_), .A2(KEYINPUT32), .A3(new_n403_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT32), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n397_), .B1(new_n425_), .B2(new_n402_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n373_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT94), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n373_), .A2(new_n426_), .A3(new_n424_), .A4(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n369_), .B(KEYINPUT33), .ZN(new_n431_));
  INV_X1    g230(.A(new_n353_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n361_), .A2(new_n432_), .A3(new_n362_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n352_), .B(new_n433_), .C1(new_n368_), .C2(new_n432_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n431_), .A2(new_n404_), .A3(new_n405_), .A4(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n428_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n375_), .A2(new_n422_), .B1(new_n423_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G232gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G29gat), .B(G36gat), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(G43gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(G43gat), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n442_), .A2(G50gat), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(G50gat), .B1(new_n442_), .B2(new_n443_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G85gat), .B(G92gat), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT9), .ZN(new_n449_));
  AND3_X1   g248(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n449_), .B(new_n452_), .C1(KEYINPUT9), .C2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT10), .B(G99gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT64), .B(G106gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT66), .B1(new_n450_), .B2(new_n451_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT66), .ZN(new_n468_));
  NAND3_X1  g267(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n464_), .A3(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n471_), .A2(KEYINPUT67), .A3(new_n448_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT67), .B1(new_n471_), .B2(new_n448_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n463_), .A2(new_n452_), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT65), .B(KEYINPUT8), .Z(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n448_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n447_), .B(new_n459_), .C1(new_n475_), .C2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n446_), .A2(KEYINPUT15), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n471_), .A2(new_n448_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n471_), .A2(KEYINPUT67), .A3(new_n448_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT8), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n458_), .B1(new_n489_), .B2(new_n478_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n480_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n491_), .A2(KEYINPUT70), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n491_), .B2(KEYINPUT70), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n440_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n490_), .A2(new_n484_), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n458_), .B(new_n446_), .C1(new_n489_), .C2(new_n478_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT70), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT34), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n491_), .A2(KEYINPUT70), .A3(new_n492_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n439_), .A3(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n495_), .A2(new_n501_), .A3(KEYINPUT35), .ZN(new_n502_));
  INV_X1    g301(.A(new_n491_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n503_), .A2(KEYINPUT35), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n438_), .B1(new_n502_), .B2(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n493_), .A2(new_n494_), .A3(new_n440_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n439_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n504_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n495_), .A2(new_n501_), .A3(KEYINPUT35), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(KEYINPUT72), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G190gat), .B(G218gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G134gat), .ZN(new_n514_));
  INV_X1    g313(.A(G162gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT71), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n507_), .A2(new_n512_), .A3(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n510_), .A2(new_n517_), .A3(new_n516_), .A4(new_n511_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT37), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n502_), .B2(new_n506_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n525_), .A3(KEYINPUT37), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT16), .B(G183gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G211gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G127gat), .B(G155gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n531_), .A2(KEYINPUT17), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT73), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536_));
  INV_X1    g335(.A(G1gat), .ZN(new_n537_));
  INV_X1    g336(.A(G8gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT14), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G8gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n535_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n544_), .A2(KEYINPUT11), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(KEYINPUT11), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G71gat), .B(G78gat), .ZN(new_n547_));
  OR3_X1    g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n547_), .A3(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n543_), .A2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n531_), .A2(KEYINPUT17), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n543_), .A2(new_n551_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n437_), .A2(new_n527_), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n490_), .B(new_n551_), .ZN(new_n558_));
  INV_X1    g357(.A(G230gat), .ZN(new_n559_));
  INV_X1    g358(.A(G233gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n287_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT5), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n206_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n490_), .A2(new_n550_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n490_), .A2(new_n550_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(KEYINPUT12), .A3(new_n570_), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n490_), .A2(KEYINPUT12), .A3(new_n550_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n564_), .B(new_n568_), .C1(new_n573_), .C2(new_n561_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n575_));
  INV_X1    g374(.A(new_n568_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n561_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n563_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT68), .B(new_n576_), .C1(new_n577_), .C2(new_n563_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT13), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(KEYINPUT13), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n542_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n446_), .A2(new_n587_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(KEYINPUT75), .B2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(KEYINPUT75), .B2(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n446_), .B(new_n587_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT74), .Z(new_n595_));
  INV_X1    g394(.A(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G169gat), .B(G197gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT76), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n231_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n579_), .A2(KEYINPUT69), .A3(new_n607_), .A4(new_n580_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n586_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n557_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n537_), .A3(new_n373_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT38), .ZN(new_n613_));
  INV_X1    g412(.A(new_n522_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n437_), .A2(new_n556_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n586_), .A2(KEYINPUT97), .A3(new_n606_), .A4(new_n608_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT98), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(new_n373_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n613_), .B1(new_n622_), .B2(new_n537_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(new_n407_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n419_), .A2(new_n420_), .A3(new_n416_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n420_), .B1(new_n419_), .B2(new_n416_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n611_), .A2(new_n538_), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G8gat), .B1(new_n620_), .B2(new_n422_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(KEYINPUT39), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n611_), .A2(new_n638_), .A3(new_n255_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n621_), .A2(new_n255_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n640_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(new_n640_), .B2(G15gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n639_), .B1(new_n641_), .B2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n335_), .A2(new_n336_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT100), .Z(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n611_), .A2(new_n644_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n621_), .A2(new_n647_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(G22gat), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT42), .B(new_n644_), .C1(new_n621_), .C2(new_n647_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(G1327gat));
  NAND2_X1  g452(.A1(new_n436_), .A2(new_n423_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n337_), .A2(new_n348_), .A3(new_n374_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n629_), .B2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(new_n614_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n610_), .A3(new_n556_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n373_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n555_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n619_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n656_), .A2(new_n527_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n656_), .B2(new_n527_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n661_), .A2(new_n662_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n526_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n437_), .B2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n656_), .A2(new_n527_), .A3(new_n666_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n670_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n665_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n671_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(G29gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n660_), .B1(new_n680_), .B2(new_n373_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT102), .ZN(G1328gat));
  AOI21_X1  g481(.A(new_n422_), .B1(new_n671_), .B2(new_n678_), .ZN(new_n683_));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT103), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n677_), .B1(new_n676_), .B2(new_n665_), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n670_), .B(new_n664_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n629_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(G36gat), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT46), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n658_), .A2(G36gat), .A3(new_n422_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n685_), .A2(new_n690_), .A3(new_n692_), .A4(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1329gat));
  NAND3_X1  g497(.A1(new_n679_), .A2(G43gat), .A3(new_n255_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n679_), .A2(KEYINPUT107), .A3(G43gat), .A4(new_n255_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT108), .B(G43gat), .Z(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n658_), .B2(new_n347_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n702_), .A3(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g505(.A1(new_n658_), .A2(G50gat), .A3(new_n646_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n645_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n679_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n709_), .B2(G50gat), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT109), .Z(G1331gat));
  NAND2_X1  g510(.A1(new_n586_), .A2(new_n608_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n606_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n615_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n374_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n557_), .A2(new_n373_), .A3(new_n714_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(new_n718_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n715_), .B2(new_n422_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT48), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n557_), .A2(new_n714_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n422_), .A2(G64gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n715_), .B2(new_n347_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT49), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n722_), .A2(G71gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n347_), .B2(new_n727_), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n715_), .B2(new_n646_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n646_), .A2(G78gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT110), .Z(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n722_), .B2(new_n732_), .ZN(G1335gat));
  OR2_X1    g532(.A1(new_n676_), .A2(KEYINPUT112), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n713_), .A2(new_n606_), .A3(new_n555_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n676_), .A2(KEYINPUT112), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G85gat), .ZN(new_n738_));
  OR3_X1    g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n374_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n657_), .A2(new_n735_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT111), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n373_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n738_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n739_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n739_), .A2(KEYINPUT113), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1336gat));
  AOI21_X1  g547(.A(G92gat), .B1(new_n741_), .B2(new_n629_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n737_), .A2(new_n422_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g550(.A(G99gat), .B1(new_n737_), .B2(new_n347_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n741_), .A2(new_n455_), .A3(new_n255_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g554(.A1(new_n676_), .A2(new_n708_), .A3(new_n735_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n676_), .A2(KEYINPUT114), .A3(new_n708_), .A4(new_n735_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(G106gat), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT52), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n758_), .A2(new_n762_), .A3(G106gat), .A4(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n741_), .A2(new_n456_), .A3(new_n708_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n768_), .A3(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1339gat));
  INV_X1    g569(.A(new_n606_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n586_), .A2(new_n771_), .A3(new_n608_), .A4(new_n555_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n673_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT54), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n573_), .A2(new_n561_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n577_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n577_), .A2(new_n777_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n576_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n606_), .A2(KEYINPUT116), .A3(new_n574_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT116), .B1(new_n606_), .B2(new_n574_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n783_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n602_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n595_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n596_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n605_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n581_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT57), .B(new_n522_), .C1(new_n787_), .C2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n783_), .B2(new_n786_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n614_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n791_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n781_), .A2(new_n782_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n780_), .B2(new_n576_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n574_), .B(new_n798_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n673_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n556_), .B1(new_n797_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n708_), .B1(new_n775_), .B2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n629_), .A2(new_n374_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n255_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n606_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n808_), .A2(KEYINPUT59), .A3(new_n255_), .A4(new_n809_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n606_), .A2(G113gat), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT118), .Z(new_n818_));
  AOI21_X1  g617(.A(new_n812_), .B1(new_n816_), .B2(new_n818_), .ZN(G1340gat));
  OAI21_X1  g618(.A(new_n238_), .B1(new_n713_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n811_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n238_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n713_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n238_), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n811_), .B2(new_n555_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT119), .B(G127gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n555_), .A2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT120), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n816_), .B2(new_n827_), .ZN(G1342gat));
  AOI21_X1  g627(.A(G134gat), .B1(new_n811_), .B2(new_n614_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n673_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n775_), .A2(new_n807_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n645_), .A2(new_n255_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n809_), .A2(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT121), .Z(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n606_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n712_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g640(.A1(new_n836_), .A2(new_n556_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT61), .B(G155gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  NOR3_X1   g643(.A1(new_n836_), .A2(new_n515_), .A3(new_n673_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n837_), .A2(new_n614_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n515_), .B2(new_n846_), .ZN(G1347gat));
  AOI21_X1  g646(.A(new_n647_), .B1(new_n775_), .B2(new_n807_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n422_), .A2(new_n373_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n255_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n606_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G169gat), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n855_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n852_), .A2(G169gat), .A3(new_n857_), .A4(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n856_), .B(new_n859_), .C1(new_n384_), .C2(new_n852_), .ZN(G1348gat));
  NAND2_X1  g659(.A1(new_n848_), .A2(new_n851_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n206_), .A3(new_n712_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n808_), .A2(new_n712_), .A3(new_n851_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n206_), .B2(new_n864_), .ZN(G1349gat));
  NOR3_X1   g664(.A1(new_n861_), .A2(new_n209_), .A3(new_n556_), .ZN(new_n866_));
  INV_X1    g665(.A(G183gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n808_), .A2(new_n555_), .A3(new_n851_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1350gat));
  NAND3_X1  g668(.A1(new_n862_), .A2(new_n210_), .A3(new_n614_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G190gat), .B1(new_n861_), .B2(new_n673_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1351gat));
  AND3_X1   g671(.A1(new_n832_), .A2(new_n833_), .A3(new_n849_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n606_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n289_), .A2(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n289_), .A2(KEYINPUT123), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n874_), .B2(new_n876_), .ZN(G1352gat));
  NAND3_X1  g677(.A1(new_n832_), .A2(new_n833_), .A3(new_n849_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n713_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n287_), .ZN(G1353gat));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n882_));
  INV_X1    g681(.A(G211gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n555_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT124), .Z(new_n885_));
  NAND2_X1  g684(.A1(new_n873_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n882_), .A2(new_n883_), .A3(KEYINPUT125), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n889_), .B2(new_n886_), .ZN(G1354gat));
  INV_X1    g690(.A(G218gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n873_), .B2(new_n527_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n879_), .A2(G218gat), .A3(new_n522_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT126), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n873_), .A2(new_n892_), .A3(new_n614_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  OAI21_X1  g696(.A(G218gat), .B1(new_n879_), .B2(new_n673_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n899_), .ZN(G1355gat));
endmodule


