//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n980_, new_n982_, new_n983_, new_n985_,
    new_n986_, new_n988_, new_n989_, new_n990_, new_n991_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT65), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT65), .B1(new_n205_), .B2(new_n207_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n211_), .A2(KEYINPUT64), .A3(new_n212_), .A4(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G85gat), .A3(G92gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G85gat), .B(G92gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(new_n219_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n210_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n221_), .A2(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(KEYINPUT66), .A3(new_n230_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n228_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n226_), .B1(new_n210_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n205_), .A2(new_n207_), .ZN(new_n238_));
  NOR4_X1   g037(.A1(new_n232_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT66), .B1(new_n229_), .B2(new_n230_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n238_), .B(new_n227_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n221_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n237_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n224_), .B1(new_n236_), .B2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G29gat), .B(G36gat), .Z(new_n245_));
  XOR2_X1   g044(.A(G43gat), .B(G50gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G29gat), .B(G36gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G43gat), .B(G50gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n247_), .A2(KEYINPUT15), .A3(new_n250_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n244_), .A2(new_n255_), .A3(KEYINPUT71), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT71), .B1(new_n244_), .B2(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n203_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT34), .Z(new_n260_));
  INV_X1    g059(.A(KEYINPUT35), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT72), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n239_), .A2(new_n240_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n206_), .B1(G99gat), .B2(G106gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n227_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n242_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT8), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n238_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT65), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n227_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n225_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n222_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n269_), .A2(new_n275_), .B1(new_n218_), .B2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n263_), .B1(new_n277_), .B2(new_n251_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n260_), .A2(new_n261_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n258_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  OAI221_X1 g081(.A(new_n278_), .B1(new_n203_), .B2(new_n282_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G190gat), .B(G218gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G134gat), .B(G162gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT36), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT74), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n281_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n286_), .B(KEYINPUT36), .Z(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT37), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n202_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n281_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  AOI211_X1 g097(.A(KEYINPUT75), .B(new_n291_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT37), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n202_), .B(KEYINPUT37), .C1(new_n298_), .C2(new_n299_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT77), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(new_n305_), .A3(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G15gat), .B(G22gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G1gat), .A2(G8gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT14), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n308_), .A2(new_n310_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n308_), .A2(new_n309_), .A3(new_n313_), .A4(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G231gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G57gat), .B(G64gat), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(KEYINPUT11), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(KEYINPUT11), .ZN(new_n322_));
  XOR2_X1   g121(.A(G71gat), .B(G78gat), .Z(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n319_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n319_), .A2(new_n327_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT67), .B1(new_n328_), .B2(new_n329_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G183gat), .B(G211gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT79), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT80), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n336_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G155gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT17), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(KEYINPUT17), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT81), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n334_), .A2(KEYINPUT82), .A3(new_n343_), .A4(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n345_), .B(new_n343_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n330_), .B1(KEYINPUT17), .B2(new_n341_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(KEYINPUT17), .B2(new_n341_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n307_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G120gat), .B(G148gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(G176gat), .B(G204gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n244_), .A2(new_n331_), .A3(KEYINPUT12), .A4(new_n326_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT12), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n362_), .B(new_n224_), .C1(new_n236_), .C2(new_n243_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n327_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n331_), .A2(KEYINPUT12), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n269_), .A2(new_n275_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(new_n224_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n361_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G230gat), .A2(G233gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n277_), .A2(new_n327_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n369_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n244_), .A2(new_n326_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n360_), .B1(new_n370_), .B2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n327_), .B(new_n363_), .C1(new_n277_), .C2(new_n365_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n372_), .B1(new_n377_), .B2(new_n361_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n378_), .A2(new_n374_), .A3(new_n359_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT69), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n375_), .A3(new_n360_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n359_), .B1(new_n378_), .B2(new_n374_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT13), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n380_), .A2(KEYINPUT13), .A3(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT70), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n390_), .A2(KEYINPUT70), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G15gat), .B(G43gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G99gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n395_), .B(KEYINPUT90), .ZN(new_n399_));
  INV_X1    g198(.A(G99gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G71gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n402_), .B(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT24), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT25), .B(G183gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT26), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n421_), .B(G190gat), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(G190gat), .ZN(new_n425_));
  INV_X1    g224(.A(G190gat), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT85), .B(KEYINPUT26), .C1(new_n426_), .C2(KEYINPUT86), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n420_), .A2(new_n424_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n408_), .A2(new_n411_), .A3(KEYINPUT87), .A4(new_n412_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n415_), .A2(new_n419_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT88), .B(G176gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT22), .B(G169gat), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n431_), .A2(new_n432_), .B1(G169gat), .B2(G176gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n411_), .B(new_n412_), .C1(G183gat), .C2(G190gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT89), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n409_), .B(KEYINPUT23), .ZN(new_n436_));
  INV_X1    g235(.A(G183gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT89), .B1(new_n437_), .B2(new_n426_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n433_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n430_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT30), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT91), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n405_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n405_), .B2(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G127gat), .B(G134gat), .Z(new_n447_));
  XOR2_X1   g246(.A(G113gat), .B(G120gat), .Z(new_n448_));
  XOR2_X1   g247(.A(new_n447_), .B(new_n448_), .Z(new_n449_));
  NAND2_X1  g248(.A1(new_n405_), .A2(new_n442_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT92), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n405_), .A2(new_n442_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n446_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n449_), .B1(new_n446_), .B2(new_n454_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n394_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n446_), .A2(new_n454_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n447_), .B(new_n448_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n446_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n393_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G57gat), .B(G85gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT101), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(new_n311_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n467_));
  INV_X1    g266(.A(G29gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n466_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G141gat), .A2(G148gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G141gat), .A2(G148gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT94), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G155gat), .A3(G162gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G155gat), .ZN(new_n482_));
  INV_X1    g281(.A(G162gat), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n481_), .A2(KEYINPUT1), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT1), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n478_), .A2(new_n480_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n476_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n474_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT2), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n472_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n489_), .A2(new_n491_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n482_), .A2(new_n483_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n481_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n449_), .B1(new_n487_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n481_), .A2(KEYINPUT1), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n499_), .A2(new_n486_), .A3(new_n495_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n459_), .B(new_n496_), .C1(new_n500_), .C2(new_n476_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n501_), .A3(KEYINPUT4), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT99), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n496_), .B1(new_n500_), .B2(new_n476_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n449_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n502_), .A2(new_n503_), .A3(new_n505_), .A4(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n498_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n487_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n459_), .B1(new_n512_), .B2(new_n496_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n504_), .B1(new_n513_), .B2(new_n507_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n503_), .B1(new_n514_), .B2(new_n502_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n471_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n502_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n508_), .A2(new_n505_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT99), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n519_), .A2(new_n470_), .A3(new_n510_), .A4(new_n509_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT28), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n487_), .A2(new_n497_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT29), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(G197gat), .A2(G204gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G197gat), .A2(G204gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT21), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(KEYINPUT21), .A3(new_n529_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G211gat), .B(G218gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n506_), .B2(KEYINPUT29), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n524_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n527_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n543_), .B2(new_n526_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G228gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G78gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G106gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G22gat), .B(G50gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n542_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G226gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n560_));
  OR2_X1    g359(.A1(KEYINPUT88), .A2(G176gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(KEYINPUT88), .A2(G176gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n432_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n417_), .A3(new_n434_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(G190gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n420_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n416_), .A2(new_n417_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n407_), .A2(KEYINPUT96), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT24), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n566_), .B1(new_n567_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n406_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n436_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n564_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n560_), .B1(new_n575_), .B2(new_n537_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n538_), .A2(new_n430_), .A3(new_n440_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n559_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G8gat), .B(G36gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G64gat), .B(G92gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n441_), .A2(new_n537_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n418_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n566_), .A2(new_n573_), .A3(new_n436_), .A4(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n588_), .A2(new_n535_), .A3(new_n536_), .A4(new_n564_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n585_), .A2(KEYINPUT20), .A3(new_n559_), .A4(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n579_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT27), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT104), .ZN(new_n593_));
  OAI211_X1 g392(.A(KEYINPUT103), .B(KEYINPUT20), .C1(new_n575_), .C2(new_n537_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n585_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT103), .B1(new_n589_), .B2(KEYINPUT20), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n558_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n576_), .A2(new_n577_), .A3(new_n559_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n593_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT20), .B1(new_n575_), .B2(new_n537_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n585_), .A3(new_n594_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT104), .B1(new_n603_), .B2(new_n558_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n584_), .B(KEYINPUT106), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n592_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n584_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n590_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n578_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n591_), .A3(KEYINPUT98), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT27), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(new_n608_), .C1(new_n609_), .C2(new_n578_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n607_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n463_), .A2(new_n522_), .A3(new_n555_), .A4(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n554_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n607_), .A2(new_n618_), .A3(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n584_), .A2(KEYINPUT32), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n599_), .B2(new_n604_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n620_), .B(KEYINPUT102), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n579_), .A3(new_n590_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n521_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n521_), .A2(new_n622_), .A3(KEYINPUT105), .A4(new_n624_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n520_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n611_), .A2(new_n614_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n520_), .A2(new_n629_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n502_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n498_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n471_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .A4(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n627_), .A2(new_n628_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n619_), .B1(new_n637_), .B2(new_n555_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n617_), .B1(new_n638_), .B2(new_n463_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G113gat), .B(G141gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G169gat), .B(G197gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n640_), .B(new_n641_), .Z(new_n642_));
  INV_X1    g441(.A(new_n316_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n250_), .B(new_n247_), .C1(new_n643_), .C2(new_n314_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n251_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT83), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n644_), .A2(new_n645_), .A3(KEYINPUT83), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n253_), .A2(new_n317_), .A3(new_n254_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(new_n649_), .A3(new_n645_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n642_), .B1(new_n655_), .B2(KEYINPUT84), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT84), .ZN(new_n657_));
  INV_X1    g456(.A(new_n642_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n657_), .B(new_n658_), .C1(new_n652_), .C2(new_n654_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n639_), .A2(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n354_), .A2(new_n391_), .A3(new_n392_), .A4(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n522_), .A2(G1gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT107), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n293_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n639_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n660_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n389_), .A2(new_n353_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G1gat), .B1(new_n673_), .B2(new_n522_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT108), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n665_), .A2(KEYINPUT107), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n665_), .A2(KEYINPUT107), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(KEYINPUT38), .A3(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n668_), .A2(new_n675_), .A3(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(new_n616_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n663_), .A2(new_n312_), .A3(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n670_), .A2(new_n680_), .A3(new_n672_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G8gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G8gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g486(.A(new_n463_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G15gat), .B1(new_n673_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OR3_X1    g490(.A1(new_n662_), .A2(G15gat), .A3(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n690_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(G1326gat));
  OR3_X1    g493(.A1(new_n662_), .A2(G22gat), .A3(new_n555_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G22gat), .B1(new_n673_), .B2(new_n555_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT42), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT42), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(G1327gat));
  AND3_X1   g498(.A1(new_n301_), .A2(new_n305_), .A3(new_n302_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n305_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n639_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT43), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n639_), .B(new_n704_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n390_), .A2(new_n660_), .A3(new_n353_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT44), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n710_), .B(new_n707_), .C1(new_n703_), .C2(new_n705_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n709_), .A2(new_n711_), .A3(new_n522_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n353_), .A2(new_n293_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n389_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n661_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n521_), .A2(new_n468_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT110), .ZN(new_n717_));
  OAI22_X1  g516(.A1(new_n712_), .A2(new_n468_), .B1(new_n715_), .B2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  INV_X1    g518(.A(G36gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n709_), .A2(new_n711_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n680_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n680_), .A2(KEYINPUT111), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n680_), .A2(KEYINPUT111), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n661_), .A2(new_n720_), .A3(new_n714_), .A4(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n726_), .B(new_n727_), .Z(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n719_), .B1(new_n722_), .B2(new_n729_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n709_), .A2(new_n711_), .A3(new_n616_), .ZN(new_n731_));
  OAI211_X1 g530(.A(KEYINPUT46), .B(new_n728_), .C1(new_n731_), .C2(new_n720_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1329gat));
  INV_X1    g532(.A(G43gat), .ZN(new_n734_));
  NOR4_X1   g533(.A1(new_n709_), .A2(new_n711_), .A3(new_n734_), .A4(new_n688_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n715_), .A2(new_n688_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(G43gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT47), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n688_), .A2(new_n734_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n721_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(G1330gat));
  INV_X1    g542(.A(G50gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n555_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n661_), .A2(new_n554_), .A3(new_n714_), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n721_), .A2(new_n745_), .B1(new_n744_), .B2(new_n746_), .ZN(G1331gat));
  AOI211_X1 g546(.A(new_n660_), .B(new_n353_), .C1(new_n392_), .C2(new_n391_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n521_), .A3(new_n670_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G57gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n354_), .A2(new_n389_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT113), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT113), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n639_), .A2(new_n671_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n522_), .A2(G57gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n750_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  NAND3_X1  g556(.A1(new_n748_), .A2(new_n670_), .A3(new_n725_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G64gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT48), .ZN(new_n760_));
  INV_X1    g559(.A(new_n725_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n761_), .A2(G64gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n755_), .B2(new_n762_), .ZN(G1333gat));
  NAND3_X1  g562(.A1(new_n748_), .A2(new_n463_), .A3(new_n670_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G71gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n765_), .B(new_n766_), .Z(new_n767_));
  OR2_X1    g566(.A1(new_n688_), .A2(G71gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n755_), .B2(new_n768_), .ZN(G1334gat));
  NAND3_X1  g568(.A1(new_n748_), .A2(new_n554_), .A3(new_n670_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G78gat), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT115), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(KEYINPUT50), .A3(new_n773_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n555_), .A2(G78gat), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n776_), .B(new_n777_), .C1(new_n755_), .C2(new_n778_), .ZN(G1335gat));
  AOI21_X1  g578(.A(new_n713_), .B1(new_n392_), .B2(new_n391_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n754_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(G85gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n521_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n353_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n390_), .A2(new_n785_), .A3(new_n660_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n705_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n704_), .B1(new_n307_), .B2(new_n639_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT116), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n706_), .A2(new_n791_), .A3(new_n786_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n522_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n784_), .B1(new_n793_), .B2(new_n783_), .ZN(G1336gat));
  INV_X1    g593(.A(G92gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n782_), .A2(new_n795_), .A3(new_n680_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n761_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n795_), .ZN(G1337gat));
  AOI21_X1  g597(.A(new_n688_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n463_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n800_));
  OAI22_X1  g599(.A1(new_n799_), .A2(new_n400_), .B1(new_n781_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  OAI221_X1 g603(.A(new_n802_), .B1(new_n781_), .B2(new_n800_), .C1(new_n799_), .C2(new_n400_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n706_), .A2(new_n554_), .A3(new_n786_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(new_n808_), .A3(G106gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(G106gat), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n554_), .A2(new_n212_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n809_), .A2(new_n810_), .B1(new_n781_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT53), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814_));
  OAI221_X1 g613(.A(new_n814_), .B1(new_n781_), .B2(new_n811_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT123), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n389_), .A2(new_n353_), .A3(new_n660_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n304_), .A2(new_n818_), .A3(new_n306_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n653_), .A2(new_n650_), .A3(new_n645_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  MUX2_X1   g623(.A(new_n655_), .B(new_n824_), .S(new_n658_), .Z(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n379_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT120), .B1(new_n370_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n378_), .A2(new_n831_), .A3(KEYINPUT55), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n369_), .B1(new_n368_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n377_), .A2(KEYINPUT119), .A3(new_n361_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n835_), .A2(new_n836_), .B1(new_n370_), .B2(new_n829_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n828_), .B(new_n360_), .C1(new_n833_), .C2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n370_), .A2(new_n829_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n368_), .A2(new_n834_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n836_), .A3(new_n372_), .ZN(new_n841_));
  AND4_X1   g640(.A1(new_n831_), .A2(new_n368_), .A3(KEYINPUT55), .A4(new_n369_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n831_), .B1(new_n378_), .B2(KEYINPUT55), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n839_), .B(new_n841_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n844_), .B2(new_n359_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n827_), .B1(new_n838_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n827_), .B(KEYINPUT58), .C1(new_n838_), .C2(new_n845_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n848_), .B(new_n849_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n376_), .A2(new_n379_), .A3(KEYINPUT69), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n825_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT121), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n385_), .A2(new_n855_), .A3(new_n825_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n660_), .A2(new_n381_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n660_), .A2(KEYINPUT118), .A3(new_n381_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n844_), .A2(new_n359_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n828_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n844_), .A2(KEYINPUT56), .A3(new_n359_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n669_), .B1(new_n857_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n861_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT118), .B1(new_n660_), .B2(new_n381_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n838_), .B2(new_n845_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n856_), .A3(new_n854_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(KEYINPUT57), .A3(new_n669_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n850_), .A2(new_n869_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n785_), .B1(new_n876_), .B2(KEYINPUT122), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n850_), .A2(new_n878_), .A3(new_n869_), .A4(new_n875_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n821_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n688_), .A2(new_n522_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n680_), .A2(new_n554_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n817_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n869_), .A2(new_n875_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n848_), .A2(new_n849_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(new_n353_), .A3(new_n879_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n700_), .A2(new_n701_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n820_), .A3(new_n818_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n819_), .A2(KEYINPUT54), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n883_), .B1(new_n889_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT123), .ZN(new_n895_));
  INV_X1    g694(.A(G113gat), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n884_), .A2(new_n895_), .A3(new_n896_), .A4(new_n660_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n876_), .A2(new_n353_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n893_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n883_), .A2(KEYINPUT59), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n660_), .B(new_n901_), .C1(new_n894_), .C2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n897_), .B1(new_n904_), .B2(new_n896_), .ZN(G1340gat));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT60), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n390_), .B2(KEYINPUT60), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n884_), .A2(new_n895_), .A3(new_n907_), .A4(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n392_), .A2(new_n391_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n910_), .B(new_n901_), .C1(new_n894_), .C2(new_n902_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n909_), .B1(new_n912_), .B2(new_n906_), .ZN(G1341gat));
  NAND3_X1  g712(.A1(new_n884_), .A2(new_n895_), .A3(new_n785_), .ZN(new_n914_));
  INV_X1    g713(.A(G127gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n889_), .A2(new_n893_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n883_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n918_), .A2(KEYINPUT59), .B1(new_n899_), .B2(new_n900_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n915_), .B1(new_n785_), .B2(KEYINPUT124), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(KEYINPUT124), .B2(new_n915_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n914_), .A2(new_n915_), .B1(new_n919_), .B2(new_n921_), .ZN(G1342gat));
  INV_X1    g721(.A(G134gat), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n884_), .A2(new_n895_), .A3(new_n923_), .A4(new_n293_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n307_), .B(new_n901_), .C1(new_n894_), .C2(new_n902_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n926_), .B2(new_n923_), .ZN(G1343gat));
  NOR3_X1   g726(.A1(new_n725_), .A2(new_n522_), .A3(new_n555_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n916_), .A2(new_n688_), .A3(new_n660_), .A4(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT125), .B(G141gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1344gat));
  NOR2_X1   g730(.A1(new_n880_), .A2(new_n463_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n932_), .A2(new_n910_), .A3(new_n928_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G148gat), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n916_), .A2(new_n688_), .A3(new_n928_), .ZN(new_n935_));
  INV_X1    g734(.A(G148gat), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n935_), .A2(new_n936_), .A3(new_n910_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(G1345gat));
  NAND3_X1  g737(.A1(new_n932_), .A2(new_n785_), .A3(new_n928_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n935_), .A2(new_n785_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1346gat));
  NAND2_X1  g743(.A1(new_n935_), .A2(new_n293_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n890_), .A2(new_n483_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT126), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n945_), .A2(new_n483_), .B1(new_n935_), .B2(new_n947_), .ZN(G1347gat));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n688_), .A2(new_n521_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n725_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n554_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n855_), .B1(new_n385_), .B2(new_n825_), .ZN(new_n953_));
  AOI211_X1 g752(.A(KEYINPUT121), .B(new_n826_), .C1(new_n380_), .C2(new_n384_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  AOI211_X1 g754(.A(new_n868_), .B(new_n293_), .C1(new_n955_), .C2(new_n873_), .ZN(new_n956_));
  AOI21_X1  g755(.A(KEYINPUT57), .B1(new_n874_), .B2(new_n669_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n785_), .B1(new_n958_), .B2(new_n850_), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n660_), .B(new_n952_), .C1(new_n821_), .C2(new_n959_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n960_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n961_));
  INV_X1    g760(.A(new_n952_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n898_), .B2(new_n893_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n963_), .A2(new_n432_), .A3(new_n660_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n961_), .A2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(KEYINPUT62), .B1(new_n960_), .B2(G169gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n949_), .B1(new_n965_), .B2(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n960_), .A2(G169gat), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  NAND4_X1  g769(.A1(new_n970_), .A2(KEYINPUT127), .A3(new_n964_), .A4(new_n961_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n967_), .A2(new_n971_), .ZN(G1348gat));
  NOR2_X1   g771(.A1(new_n880_), .A2(new_n554_), .ZN(new_n973_));
  INV_X1    g772(.A(new_n951_), .ZN(new_n974_));
  AND3_X1   g773(.A1(new_n974_), .A2(G176gat), .A3(new_n910_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n963_), .A2(new_n389_), .ZN(new_n976_));
  AOI22_X1  g775(.A1(new_n973_), .A2(new_n975_), .B1(new_n431_), .B2(new_n976_), .ZN(G1349gat));
  INV_X1    g776(.A(new_n963_), .ZN(new_n978_));
  NOR3_X1   g777(.A1(new_n978_), .A2(new_n420_), .A3(new_n353_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n973_), .A2(new_n785_), .A3(new_n974_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n979_), .B1(new_n980_), .B2(new_n437_), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n978_), .B2(new_n890_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n963_), .A2(new_n565_), .A3(new_n293_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n982_), .A2(new_n983_), .ZN(G1351gat));
  NOR2_X1   g783(.A1(new_n761_), .A2(new_n618_), .ZN(new_n985_));
  NAND4_X1  g784(.A1(new_n916_), .A2(new_n688_), .A3(new_n660_), .A4(new_n985_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g786(.A1(new_n932_), .A2(new_n910_), .A3(new_n985_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n988_), .A2(G204gat), .ZN(new_n989_));
  INV_X1    g788(.A(G204gat), .ZN(new_n990_));
  NAND4_X1  g789(.A1(new_n932_), .A2(new_n990_), .A3(new_n910_), .A4(new_n985_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n989_), .A2(new_n991_), .ZN(G1353gat));
  XOR2_X1   g791(.A(KEYINPUT63), .B(G211gat), .Z(new_n993_));
  NAND4_X1  g792(.A1(new_n932_), .A2(new_n785_), .A3(new_n985_), .A4(new_n993_), .ZN(new_n994_));
  NAND4_X1  g793(.A1(new_n916_), .A2(new_n688_), .A3(new_n785_), .A4(new_n985_), .ZN(new_n995_));
  NOR2_X1   g794(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n995_), .A2(new_n996_), .ZN(new_n997_));
  AND2_X1   g796(.A1(new_n994_), .A2(new_n997_), .ZN(G1354gat));
  NAND3_X1  g797(.A1(new_n932_), .A2(new_n307_), .A3(new_n985_), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n999_), .A2(G218gat), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(new_n669_), .A2(G218gat), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n932_), .A2(new_n985_), .A3(new_n1001_), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n1000_), .A2(new_n1002_), .ZN(G1355gat));
endmodule


