//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT83), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G15gat), .B(G43gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT82), .ZN(new_n206_));
  XOR2_X1   g005(.A(G71gat), .B(G99gat), .Z(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT79), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n213_), .A2(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI221_X1 g017(.A(KEYINPUT80), .B1(G183gat), .B2(G190gat), .C1(new_n213_), .C2(new_n215_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G169gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT78), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n224_), .A3(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(new_n228_), .A3(new_n221_), .A4(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n218_), .A2(new_n219_), .A3(new_n223_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n220_), .A2(new_n221_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n210_), .A2(new_n212_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n232_), .A2(KEYINPUT24), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(G183gat), .ZN(new_n240_));
  INV_X1    g039(.A(G183gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT25), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n240_), .B(new_n242_), .C1(KEYINPUT76), .C2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(KEYINPUT76), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(KEYINPUT77), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n238_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n231_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n230_), .A2(new_n223_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n257_), .A2(new_n219_), .B1(new_n238_), .B2(new_n250_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n253_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n208_), .B1(new_n260_), .B2(KEYINPUT84), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n231_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n253_), .B1(new_n231_), .B2(new_n251_), .ZN(new_n263_));
  OAI211_X1 g062(.A(KEYINPUT84), .B(new_n208_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n204_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n260_), .A2(KEYINPUT84), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT84), .B1(new_n262_), .B2(new_n263_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n208_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n203_), .A3(new_n264_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(new_n267_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT86), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G113gat), .B(G120gat), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n275_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(KEYINPUT85), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT85), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n275_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT31), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n273_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n271_), .A2(new_n267_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n203_), .B1(new_n270_), .B2(new_n264_), .ZN(new_n286_));
  OAI211_X1 g085(.A(KEYINPUT86), .B(new_n282_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT100), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n241_), .A2(KEYINPUT25), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n239_), .A2(G183gat), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT93), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT93), .B1(new_n290_), .B2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n246_), .A2(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n244_), .A2(new_n294_), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n292_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT94), .B1(new_n296_), .B2(new_n234_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT93), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n244_), .A2(new_n294_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT93), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT94), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n233_), .ZN(new_n304_));
  OAI22_X1  g103(.A1(new_n213_), .A2(new_n215_), .B1(KEYINPUT24), .B2(new_n232_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n297_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT95), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n224_), .A2(G169gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n225_), .A2(new_n229_), .A3(KEYINPUT95), .ZN(new_n312_));
  AOI21_X1  g111(.A(G176gat), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT96), .B1(new_n313_), .B2(new_n222_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n236_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n225_), .A2(new_n229_), .A3(KEYINPUT95), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT95), .B1(new_n225_), .B2(new_n229_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n221_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT96), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n223_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n307_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n329_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n327_), .A2(new_n330_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n328_), .A2(new_n329_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n326_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n323_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n231_), .A3(new_n251_), .ZN(new_n343_));
  AND4_X1   g142(.A1(KEYINPUT20), .A2(new_n339_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n307_), .A2(new_n337_), .A3(new_n322_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT20), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT99), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT99), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n348_), .A3(KEYINPUT20), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n252_), .A2(new_n338_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n344_), .B1(new_n351_), .B2(new_n341_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G8gat), .B(G36gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n289_), .B1(new_n352_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n357_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n346_), .A2(KEYINPUT99), .B1(new_n338_), .B2(new_n252_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n342_), .B1(new_n360_), .B2(new_n349_), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT100), .B(new_n359_), .C1(new_n361_), .C2(new_n344_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n311_), .A2(new_n312_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n222_), .B1(new_n363_), .B2(new_n221_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n315_), .B1(new_n364_), .B2(new_n320_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n302_), .A2(new_n233_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n305_), .B1(new_n366_), .B2(KEYINPUT94), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n314_), .A2(new_n365_), .B1(new_n367_), .B2(new_n304_), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT20), .B(new_n343_), .C1(new_n368_), .C2(new_n337_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n341_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n350_), .A2(KEYINPUT20), .A3(new_n345_), .A4(new_n342_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n357_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT27), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n358_), .A2(new_n362_), .A3(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G155gat), .B(G162gat), .Z(new_n376_));
  NOR2_X1   g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT88), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT88), .ZN(new_n380_));
  OAI22_X1  g179(.A1(new_n380_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n381_));
  INV_X1    g180(.A(G141gat), .ZN(new_n382_));
  INV_X1    g181(.A(G148gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n379_), .B(new_n381_), .C1(KEYINPUT2), .C2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT89), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n376_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n384_), .B1(KEYINPUT87), .B2(new_n377_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n377_), .A2(KEYINPUT87), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n281_), .A2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n276_), .A2(new_n277_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT4), .B1(new_n396_), .B2(new_n398_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n281_), .A2(new_n395_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n400_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G85gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT0), .B(G57gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n401_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n337_), .B1(KEYINPUT29), .B2(new_n395_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G22gat), .B(G50gat), .Z(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n416_), .A2(new_n417_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n419_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n417_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n388_), .A2(new_n394_), .A3(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT28), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(KEYINPUT28), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT90), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n432_), .A3(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(G78gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n439_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n431_), .A2(new_n441_), .A3(new_n433_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n425_), .A2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n420_), .A2(new_n440_), .A3(new_n424_), .A4(new_n442_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n415_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n323_), .B2(new_n338_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n342_), .B1(new_n448_), .B2(new_n343_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n342_), .B1(new_n258_), .B2(new_n337_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n346_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n359_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n372_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT27), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT101), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT101), .ZN(new_n456_));
  AOI211_X1 g255(.A(new_n456_), .B(KEYINPUT27), .C1(new_n452_), .C2(new_n372_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n375_), .B(new_n446_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n399_), .A2(new_n400_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n411_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n400_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT33), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n413_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n407_), .A2(KEYINPUT33), .A3(new_n412_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n372_), .A3(new_n452_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n357_), .A2(KEYINPUT32), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n370_), .A2(new_n371_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT98), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n370_), .A2(new_n469_), .A3(new_n371_), .A4(new_n466_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n415_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n352_), .A2(new_n466_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n465_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n444_), .A2(new_n445_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n288_), .B1(new_n458_), .B2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n375_), .B(new_n475_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n415_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n287_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n282_), .B1(new_n272_), .B2(KEYINPUT86), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G29gat), .B(G36gat), .Z(new_n485_));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT15), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  INV_X1    g288(.A(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G8gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n487_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(new_n495_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n499_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT75), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT74), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n504_), .B(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n484_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513_));
  INV_X1    g312(.A(G85gat), .ZN(new_n514_));
  INV_X1    g313(.A(G92gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524_));
  INV_X1    g323(.A(G99gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n438_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n523_), .B1(new_n528_), .B2(KEYINPUT66), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(KEYINPUT66), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n520_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n528_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n521_), .B(KEYINPUT6), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n518_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT65), .B(G106gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT10), .B(G99gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT64), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(KEYINPUT64), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n536_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n516_), .A2(KEYINPUT9), .A3(new_n517_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n517_), .A2(KEYINPUT9), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  OAI22_X1  g345(.A1(new_n535_), .A2(KEYINPUT8), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n488_), .B1(new_n532_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT66), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n534_), .B1(new_n533_), .B2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT8), .B(new_n519_), .C1(new_n550_), .C2(new_n530_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n543_), .A2(new_n546_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n519_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT8), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n551_), .A2(new_n552_), .A3(new_n487_), .A4(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT34), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT35), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT70), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n548_), .A2(new_n556_), .A3(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n559_), .A2(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G190gat), .B(G218gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT69), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n563_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n548_), .A2(new_n569_), .A3(new_n556_), .A4(new_n561_), .ZN(new_n570_));
  AND4_X1   g369(.A1(new_n513_), .A2(new_n564_), .A3(new_n568_), .A4(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n568_), .B(new_n513_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT37), .B1(new_n574_), .B2(KEYINPUT71), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  NOR4_X1   g376(.A1(new_n571_), .A2(new_n573_), .A3(new_n576_), .A4(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n583_));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n495_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT17), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n595_), .A2(KEYINPUT17), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n590_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT73), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  NAND4_X1  g405(.A1(new_n551_), .A2(new_n552_), .A3(new_n555_), .A4(new_n587_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n585_), .A2(new_n586_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n547_), .B2(new_n532_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n609_), .A3(KEYINPUT12), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n608_), .B(new_n611_), .C1(new_n547_), .C2(new_n532_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n610_), .A2(new_n612_), .B1(G230gat), .B2(G233gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n606_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n612_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n617_), .B2(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n606_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT67), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT67), .ZN(new_n621_));
  NOR4_X1   g420(.A1(new_n613_), .A2(new_n621_), .A3(new_n615_), .A4(new_n606_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n616_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT68), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n628_));
  OAI221_X1 g427(.A(new_n616_), .B1(new_n628_), .B2(new_n625_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n580_), .A2(new_n602_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n512_), .A2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(G1gat), .A3(new_n479_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT38), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n351_), .A2(new_n341_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n344_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n357_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n373_), .B1(new_n638_), .B2(KEYINPUT100), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n449_), .A2(new_n451_), .A3(new_n359_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n357_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n454_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n456_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n453_), .A2(KEYINPUT101), .A3(new_n454_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n358_), .A2(new_n639_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n645_), .A2(new_n479_), .A3(new_n475_), .A4(new_n288_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n466_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n361_), .B2(new_n344_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(new_n415_), .A3(new_n470_), .A4(new_n468_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n474_), .B1(new_n649_), .B2(new_n465_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n645_), .B2(new_n446_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n646_), .B1(new_n651_), .B2(new_n288_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n574_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n511_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n600_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n654_), .B2(new_n600_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n653_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n479_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n634_), .A2(new_n635_), .A3(new_n660_), .ZN(G1324gat));
  XNOR2_X1  g460(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n664_), .B(G8gat), .C1(new_n659_), .C2(new_n645_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n484_), .A2(new_n574_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n645_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n658_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n670_), .A2(KEYINPUT104), .A3(new_n664_), .A4(G8gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n667_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G8gat), .B1(new_n659_), .B2(new_n645_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(KEYINPUT103), .A3(KEYINPUT39), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT103), .B1(new_n673_), .B2(KEYINPUT39), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n672_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n632_), .A2(G8gat), .A3(new_n645_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n663_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n677_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n674_), .A2(new_n675_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n679_), .B(new_n662_), .C1(new_n680_), .C2(new_n672_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1325gat));
  INV_X1    g481(.A(new_n288_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G15gat), .B1(new_n659_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n685_), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n632_), .A2(G15gat), .A3(new_n683_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(G1326gat));
  OR3_X1    g488(.A1(new_n632_), .A2(G22gat), .A3(new_n475_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G22gat), .B1(new_n659_), .B2(new_n475_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT42), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n691_), .A2(KEYINPUT42), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT107), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n697_), .B(new_n690_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1327gat));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n602_), .A2(new_n654_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n580_), .B1(new_n477_), .B2(new_n483_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n579_), .B2(KEYINPUT108), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n580_), .B(new_n703_), .C1(new_n477_), .C2(new_n483_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n700_), .B(new_n701_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n415_), .A2(G29gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n701_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n703_), .B1(new_n652_), .B2(new_n580_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n706_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(KEYINPUT109), .A3(new_n700_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(KEYINPUT44), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n707_), .B(new_n708_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n630_), .A2(new_n601_), .A3(new_n653_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n512_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G29gat), .B1(new_n720_), .B2(new_n415_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n717_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723_));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n713_), .A2(new_n716_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n715_), .A2(KEYINPUT44), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n723_), .B(new_n724_), .C1(new_n727_), .C2(new_n708_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n722_), .A2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n707_), .A2(new_n645_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n725_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n669_), .A2(new_n731_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n719_), .A2(KEYINPUT45), .A3(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT45), .B1(new_n719_), .B2(new_n734_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n730_), .B1(new_n733_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n726_), .A2(new_n669_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n716_), .B2(new_n713_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT46), .B(new_n737_), .C1(new_n741_), .C2(new_n731_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1329gat));
  NAND2_X1  g542(.A1(new_n288_), .A2(G43gat), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n707_), .B(new_n744_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G43gat), .B1(new_n720_), .B2(new_n288_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT47), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  INV_X1    g547(.A(new_n746_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n748_), .B(new_n749_), .C1(new_n727_), .C2(new_n744_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n720_), .B2(new_n474_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n727_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n474_), .A2(G50gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(G1331gat));
  NAND2_X1  g554(.A1(new_n630_), .A2(new_n511_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n668_), .A2(new_n601_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n415_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G57gat), .ZN(new_n763_));
  INV_X1    g562(.A(new_n511_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n484_), .A2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(new_n630_), .A3(new_n579_), .A4(new_n601_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n479_), .A2(G57gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1332gat));
  OR3_X1    g567(.A1(new_n766_), .A2(G64gat), .A3(new_n645_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n669_), .A3(new_n761_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(G64gat), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G64gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1333gat));
  OR3_X1    g573(.A1(new_n766_), .A2(G71gat), .A3(new_n683_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n760_), .A2(new_n288_), .A3(new_n761_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G71gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G71gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1334gat));
  NAND3_X1  g579(.A1(new_n760_), .A2(new_n474_), .A3(new_n761_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G78gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G78gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n474_), .A2(new_n436_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n783_), .A2(new_n784_), .B1(new_n766_), .B2(new_n785_), .ZN(G1335gat));
  NAND2_X1  g585(.A1(new_n757_), .A2(new_n602_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n514_), .B1(new_n788_), .B2(new_n415_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n602_), .A2(new_n630_), .A3(new_n574_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n765_), .A2(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n792_), .A2(G85gat), .A3(new_n479_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT113), .Z(G1336gat));
  AND2_X1   g594(.A1(new_n788_), .A2(new_n669_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n669_), .A2(new_n515_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n796_), .A2(new_n515_), .B1(new_n792_), .B2(new_n797_), .ZN(G1337gat));
  AND2_X1   g597(.A1(new_n539_), .A2(new_n542_), .ZN(new_n799_));
  OR3_X1    g598(.A1(new_n792_), .A2(new_n683_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n788_), .A2(new_n288_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n801_), .B2(G99gat), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n525_), .C1(new_n788_), .C2(new_n288_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT115), .A3(KEYINPUT51), .ZN(new_n806_));
  NAND2_X1  g605(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n800_), .C1(new_n802_), .C2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1338gat));
  AOI21_X1  g608(.A(new_n438_), .B1(new_n788_), .B2(new_n474_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n810_), .A2(KEYINPUT52), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(KEYINPUT52), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n475_), .A2(new_n536_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n765_), .A2(new_n791_), .A3(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT116), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT53), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n811_), .A2(new_n815_), .A3(new_n818_), .A4(new_n812_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1339gat));
  INV_X1    g619(.A(new_n620_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n622_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n496_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n501_), .A2(new_n499_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  MUX2_X1   g625(.A(new_n826_), .B(new_n504_), .S(new_n509_), .Z(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n617_), .A2(new_n614_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n613_), .B2(KEYINPUT55), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n617_), .A2(new_n614_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n613_), .A2(KEYINPUT55), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .A4(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n606_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(KEYINPUT56), .A3(new_n606_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n828_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n579_), .B1(new_n841_), .B2(KEYINPUT58), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(KEYINPUT58), .B2(new_n841_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n823_), .A2(new_n764_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n623_), .A2(new_n827_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n653_), .C1(new_n845_), .C2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n843_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n653_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n849_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n631_), .B2(new_n511_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n631_), .A2(new_n857_), .A3(new_n511_), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n856_), .A2(new_n600_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n683_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n843_), .A2(new_n848_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n852_), .A2(new_n855_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n601_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n859_), .A2(new_n858_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n861_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(KEYINPUT59), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n862_), .A2(KEYINPUT59), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n511_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n600_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n764_), .B(new_n861_), .C1(new_n873_), .C2(new_n866_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n871_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(KEYINPUT120), .A3(new_n871_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n870_), .A2(new_n872_), .B1(new_n877_), .B2(new_n878_), .ZN(G1340gat));
  OAI21_X1  g678(.A(new_n869_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n863_), .A2(new_n864_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n600_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n866_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n868_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n630_), .B(new_n880_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G120gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n888_));
  AOI21_X1  g687(.A(G120gat), .B1(new_n630_), .B2(new_n888_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n888_), .A2(G120gat), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n862_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n891_), .ZN(G1341gat));
  OAI211_X1 g691(.A(new_n600_), .B(new_n880_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G127gat), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n862_), .A2(G127gat), .A3(new_n602_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1342gat));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n579_), .A2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT122), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n574_), .B(new_n861_), .C1(new_n873_), .C2(new_n866_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n897_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n900_), .A2(KEYINPUT121), .A3(new_n897_), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n870_), .A2(new_n899_), .B1(new_n903_), .B2(new_n904_), .ZN(G1343gat));
  NOR4_X1   g704(.A1(new_n669_), .A2(new_n288_), .A3(new_n479_), .A4(new_n475_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n860_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n511_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT123), .B(G141gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1344gat));
  INV_X1    g709(.A(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n630_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G148gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n383_), .A3(new_n630_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1345gat));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n860_), .A2(new_n916_), .A3(new_n601_), .A4(new_n906_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n601_), .B(new_n906_), .C1(new_n873_), .C2(new_n866_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT124), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT61), .B(G155gat), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n917_), .A2(new_n919_), .A3(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n907_), .B2(new_n579_), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n653_), .A2(G162gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n907_), .B2(new_n925_), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n645_), .A2(new_n482_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n474_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n764_), .B(new_n929_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n930_), .A2(new_n931_), .A3(G169gat), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n867_), .A2(new_n764_), .A3(new_n363_), .A4(new_n929_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n930_), .B2(G169gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1348gat));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n883_), .B2(new_n474_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n860_), .A2(KEYINPUT125), .A3(new_n475_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n927_), .A2(G176gat), .A3(new_n630_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n867_), .A2(new_n630_), .A3(new_n929_), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n939_), .A2(new_n940_), .B1(new_n221_), .B2(new_n941_), .ZN(G1349gat));
  AOI21_X1  g741(.A(new_n882_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n867_), .A2(new_n929_), .A3(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n928_), .A2(new_n602_), .ZN(new_n945_));
  AOI21_X1  g744(.A(KEYINPUT125), .B1(new_n860_), .B2(new_n475_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n883_), .A2(new_n936_), .A3(new_n474_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n944_), .B1(new_n948_), .B2(new_n241_), .ZN(G1350gat));
  NOR2_X1   g748(.A1(new_n653_), .A2(new_n295_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n867_), .A2(new_n929_), .A3(new_n950_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n580_), .B(new_n929_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(G190gat), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n951_), .A2(KEYINPUT126), .A3(new_n953_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1351gat));
  NOR3_X1   g757(.A1(new_n288_), .A2(new_n415_), .A3(new_n475_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n669_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n883_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(new_n764_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n630_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g764(.A(new_n960_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n860_), .A2(new_n600_), .A3(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n968_));
  AND2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n967_), .A2(new_n968_), .A3(new_n969_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n970_), .B1(new_n967_), .B2(new_n968_), .ZN(G1354gat));
  AND3_X1   g770(.A1(new_n961_), .A2(G218gat), .A3(new_n580_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n961_), .A2(new_n574_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(KEYINPUT127), .ZN(new_n974_));
  NOR3_X1   g773(.A1(new_n883_), .A2(new_n653_), .A3(new_n960_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976_));
  AOI21_X1  g775(.A(G218gat), .B1(new_n975_), .B2(new_n976_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n972_), .B1(new_n974_), .B2(new_n977_), .ZN(G1355gat));
endmodule


