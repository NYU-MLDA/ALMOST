//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n203_), .B1(G155gat), .B2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT77), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT1), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT77), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G141gat), .B(G148gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OR3_X1    g014(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  INV_X1    g016(.A(G141gat), .ZN(new_n218_));
  INV_X1    g017(.A(G148gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n216_), .A2(new_n220_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227_));
  INV_X1    g026(.A(G134gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G127gat), .ZN(new_n229_));
  INV_X1    g028(.A(G127gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G134gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT75), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n227_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n230_), .A2(G134gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n228_), .A2(G127gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT75), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n227_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  AND4_X1   g041(.A1(new_n202_), .A2(new_n215_), .A3(new_n226_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n215_), .A2(new_n226_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n233_), .A2(new_n234_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n247_), .B2(new_n239_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n213_), .A2(new_n214_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n202_), .B1(new_n251_), .B2(new_n242_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT85), .B(KEYINPUT4), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n202_), .A3(new_n242_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT76), .B1(new_n235_), .B2(new_n241_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n251_), .A2(new_n260_), .A3(new_n248_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n215_), .A2(new_n242_), .A3(new_n226_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT84), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n259_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n258_), .B1(new_n264_), .B2(KEYINPUT4), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n255_), .B1(new_n265_), .B2(new_n254_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G29gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G85gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G57gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n253_), .A2(new_n272_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n254_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n270_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n255_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT93), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n271_), .A2(new_n277_), .A3(KEYINPUT93), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G15gat), .B(G43gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT74), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT30), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT23), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G169gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n292_));
  OR3_X1    g091(.A1(new_n291_), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n288_), .A2(new_n290_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT73), .B1(G169gat), .B2(G176gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(KEYINPUT73), .A2(G169gat), .A3(G176gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n295_), .B1(G169gat), .B2(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301_));
  INV_X1    g100(.A(G176gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n291_), .A3(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n303_), .A3(new_n296_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n299_), .A2(new_n288_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(KEYINPUT71), .A2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT26), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(KEYINPUT71), .A3(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(G183gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT25), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G183gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n307_), .A2(new_n309_), .A3(new_n311_), .A4(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT25), .B(G183gat), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n317_), .A2(KEYINPUT72), .A3(new_n307_), .A4(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n294_), .B1(new_n305_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n286_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(G71gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n321_), .B(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n260_), .A2(new_n248_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT31), .ZN(new_n327_));
  INV_X1    g126(.A(G99gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n329_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n283_), .A2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n244_), .A2(KEYINPUT29), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT78), .B(KEYINPUT28), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT79), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(G78gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G106gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n338_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT21), .ZN(new_n345_));
  INV_X1    g144(.A(G204gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT81), .B1(new_n346_), .B2(G197gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n350_), .B2(G197gat), .ZN(new_n351_));
  INV_X1    g150(.A(G197gat), .ZN(new_n352_));
  NOR4_X1   g151(.A1(new_n348_), .A2(new_n349_), .A3(KEYINPUT81), .A4(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n345_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n352_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n345_), .B1(G197gat), .B2(G204gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n351_), .A2(new_n353_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n355_), .A2(new_n345_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n354_), .A2(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(KEYINPUT29), .B2(new_n244_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G22gat), .B(G50gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n344_), .A2(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n338_), .A2(new_n343_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n338_), .A2(new_n343_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT18), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT19), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n362_), .B2(new_n320_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383_));
  INV_X1    g182(.A(new_n347_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT80), .B(G204gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n352_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n350_), .A2(new_n387_), .A3(G197gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n388_), .A3(new_n361_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n359_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT21), .B1(new_n386_), .B2(new_n388_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n308_), .A2(G190gat), .ZN(new_n393_));
  INV_X1    g192(.A(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT26), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n311_), .A2(new_n313_), .A3(new_n393_), .A4(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n299_), .A2(new_n304_), .A3(new_n288_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n293_), .A2(new_n292_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n287_), .B(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n400_), .B2(new_n289_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n382_), .A2(new_n383_), .B1(new_n392_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n305_), .A2(new_n319_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n401_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n392_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT82), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n380_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n362_), .A2(new_n401_), .A3(new_n397_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n392_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT20), .A4(new_n380_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n377_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n383_), .B(KEYINPUT20), .C1(new_n405_), .C2(new_n392_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n392_), .A2(new_n402_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n382_), .A2(new_n383_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n379_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n411_), .A3(new_n376_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(KEYINPUT83), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n422_), .B(new_n377_), .C1(new_n408_), .C2(new_n412_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n402_), .A2(KEYINPUT89), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT89), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n397_), .A2(new_n401_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n362_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n410_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT90), .B1(new_n428_), .B2(KEYINPUT20), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n379_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n403_), .A2(new_n380_), .A3(new_n407_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n377_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(KEYINPUT27), .A3(new_n419_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT95), .B1(new_n424_), .B2(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n424_), .A2(KEYINPUT95), .A3(new_n436_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n334_), .B(new_n372_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n271_), .A2(new_n277_), .A3(KEYINPUT93), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT93), .B1(new_n271_), .B2(new_n277_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n371_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n424_), .A2(new_n436_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n376_), .A2(KEYINPUT32), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT91), .B1(new_n434_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n450_), .B(new_n447_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n408_), .A2(new_n412_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n447_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n266_), .A2(new_n270_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n276_), .B1(new_n275_), .B2(new_n255_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n446_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n271_), .A2(new_n277_), .B1(new_n453_), .B2(new_n447_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n459_), .B(KEYINPUT92), .C1(new_n449_), .C2(new_n451_), .ZN(new_n460_));
  OR2_X1    g259(.A1(KEYINPUT86), .A2(KEYINPUT33), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n271_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT86), .A2(KEYINPUT33), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n266_), .A2(new_n270_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n420_), .A2(new_n423_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n274_), .B1(new_n253_), .B2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n467_), .B(new_n259_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n276_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT88), .B1(new_n265_), .B2(new_n254_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n265_), .A2(KEYINPUT88), .A3(new_n254_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n465_), .A2(new_n466_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n458_), .A2(new_n460_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n445_), .B1(new_n477_), .B2(new_n372_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT94), .B1(new_n478_), .B2(new_n332_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT94), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n278_), .B(new_n454_), .C1(new_n449_), .C2(new_n451_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n423_), .A2(new_n420_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n446_), .A2(new_n481_), .B1(new_n482_), .B2(new_n465_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n371_), .B1(new_n483_), .B2(new_n460_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n480_), .B(new_n333_), .C1(new_n484_), .C2(new_n445_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n440_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487_));
  INV_X1    g286(.A(G1gat), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT14), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G8gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G29gat), .B(G36gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n494_), .B(new_n495_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT15), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n493_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n500_), .B1(new_n504_), .B2(new_n499_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n505_), .B(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n486_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT5), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G176gat), .B(G204gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  NAND2_X1  g313(.A1(G230gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT10), .B(G99gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(G106gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT66), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n520_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n518_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT64), .B(G85gat), .ZN(new_n531_));
  INV_X1    g330(.A(G92gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n529_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT7), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n528_), .B2(new_n522_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G85gat), .B(G92gat), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n542_), .A2(KEYINPUT8), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n539_), .B(KEYINPUT7), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n527_), .A2(new_n520_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n519_), .A2(new_n521_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n550_), .B2(new_n543_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n538_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n556_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n552_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(new_n538_), .C1(new_n545_), .C2(new_n551_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(KEYINPUT12), .A3(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT8), .B1(new_n542_), .B2(new_n544_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n550_), .A2(new_n546_), .A3(new_n543_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n565_), .A2(new_n566_), .B1(new_n537_), .B2(new_n529_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n567_), .A2(KEYINPUT12), .A3(new_n562_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n516_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n515_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n514_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n514_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT67), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT67), .ZN(new_n575_));
  NOR4_X1   g374(.A1(new_n569_), .A2(new_n575_), .A3(new_n570_), .A4(new_n514_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n571_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n564_), .A2(new_n568_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n515_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n570_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n573_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n575_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n572_), .A2(KEYINPUT67), .A3(new_n573_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT13), .A3(new_n571_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n579_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI22_X1  g394(.A1(new_n552_), .A2(new_n496_), .B1(KEYINPUT35), .B2(new_n592_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n496_), .B(KEYINPUT15), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n567_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n595_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n567_), .A2(new_n501_), .B1(new_n594_), .B2(new_n593_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n595_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n552_), .A2(new_n502_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT68), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n606_), .B(KEYINPUT36), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT69), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n596_), .A2(new_n598_), .A3(new_n595_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n601_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n609_), .A3(new_n608_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n590_), .B1(new_n610_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n493_), .B(new_n618_), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n562_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n493_), .B(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n560_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G127gat), .B(G155gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT16), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n620_), .A2(new_n623_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(KEYINPUT70), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n631_), .B(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n611_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT37), .B1(new_n635_), .B2(new_n608_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n617_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n589_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n510_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n488_), .A3(new_n283_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n643_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n635_), .A2(new_n608_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n486_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n589_), .A2(new_n509_), .A3(new_n634_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G1gat), .B1(new_n650_), .B2(new_n282_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(new_n645_), .A3(new_n651_), .ZN(G1324gat));
  NOR2_X1   g451(.A1(new_n438_), .A2(new_n437_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n641_), .A2(new_n489_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n655_));
  INV_X1    g454(.A(new_n650_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n653_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  AND4_X1   g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .A4(G8gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n489_), .B1(KEYINPUT97), .B2(KEYINPUT39), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n657_), .A2(new_n660_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n654_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n662_), .B(new_n664_), .ZN(G1325gat));
  OR3_X1    g464(.A1(new_n640_), .A2(G15gat), .A3(new_n333_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n667_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n656_), .A2(new_n332_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n673_), .B2(G15gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n672_), .A3(G15gat), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n670_), .A2(new_n671_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n668_), .A2(new_n676_), .A3(new_n669_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT100), .B1(new_n678_), .B2(new_n674_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1326gat));
  OR3_X1    g479(.A1(new_n640_), .A2(G22gat), .A3(new_n372_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G22gat), .B1(new_n650_), .B2(new_n372_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT102), .Z(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n681_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n634_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n589_), .A2(new_n688_), .A3(new_n646_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n510_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n283_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n479_), .A2(new_n485_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n439_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n617_), .A2(new_n636_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n486_), .B2(new_n695_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n509_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n588_), .A2(new_n700_), .A3(new_n634_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT103), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT44), .B1(new_n699_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n702_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n283_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n691_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n690_), .A2(new_n710_), .A3(new_n653_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n653_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n704_), .A2(new_n706_), .A3(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n710_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n713_), .B(KEYINPUT46), .C1(new_n715_), .C2(new_n710_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1329gat));
  AOI21_X1  g519(.A(G43gat), .B1(new_n690_), .B2(new_n332_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n724_));
  INV_X1    g523(.A(G43gat), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n333_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n707_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n726_), .ZN(new_n728_));
  NOR4_X1   g527(.A1(new_n704_), .A2(new_n706_), .A3(KEYINPUT105), .A4(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n723_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT47), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(new_n723_), .C1(new_n727_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1330gat));
  NOR2_X1   g533(.A1(new_n372_), .A2(G50gat), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT108), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n690_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n707_), .A2(new_n371_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n738_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT107), .B1(new_n738_), .B2(G50gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(G1331gat));
  NAND2_X1  g540(.A1(new_n589_), .A2(new_n637_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT109), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n743_), .A2(new_n486_), .A3(new_n700_), .ZN(new_n744_));
  INV_X1    g543(.A(G57gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n283_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n648_), .A2(new_n509_), .A3(new_n589_), .A4(new_n688_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT110), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n283_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g549(.A(G64gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n744_), .A2(new_n751_), .A3(new_n653_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n748_), .A2(new_n653_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(G64gat), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT48), .B(new_n751_), .C1(new_n748_), .C2(new_n653_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1333gat));
  NAND3_X1  g556(.A1(new_n744_), .A2(new_n323_), .A3(new_n332_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n748_), .A2(new_n332_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G71gat), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT49), .B(new_n323_), .C1(new_n748_), .C2(new_n332_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(G1334gat));
  NAND3_X1  g562(.A1(new_n744_), .A2(new_n340_), .A3(new_n371_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n748_), .A2(new_n371_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G78gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT50), .B(new_n340_), .C1(new_n748_), .C2(new_n371_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n486_), .A2(new_n700_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n588_), .A2(new_n688_), .A3(new_n646_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n283_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n588_), .A2(new_n700_), .A3(new_n688_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n699_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n282_), .A2(new_n531_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT111), .Z(new_n778_));
  AOI21_X1  g577(.A(new_n774_), .B1(new_n776_), .B2(new_n778_), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n532_), .A3(new_n653_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n776_), .A2(new_n653_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n532_), .ZN(G1337gat));
  NOR3_X1   g581(.A1(new_n772_), .A2(new_n333_), .A3(new_n517_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n776_), .A2(new_n332_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(G99gat), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n773_), .A2(new_n342_), .A3(new_n371_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n699_), .A2(new_n371_), .A3(new_n775_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G106gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n564_), .A2(new_n568_), .A3(new_n516_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n581_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n580_), .A2(KEYINPUT55), .A3(new_n515_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n569_), .A2(KEYINPUT114), .A3(KEYINPUT55), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n514_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n514_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT117), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n514_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT117), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n508_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n505_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n508_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT115), .Z(new_n814_));
  AOI21_X1  g613(.A(new_n498_), .B1(new_n504_), .B2(KEYINPUT116), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(KEYINPUT116), .B2(new_n504_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n812_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n586_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n810_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n796_), .B1(new_n807_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n808_), .A2(new_n809_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n514_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n824_), .A2(KEYINPUT58), .A3(new_n810_), .A4(new_n818_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n820_), .A2(new_n696_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n509_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n577_), .A2(new_n817_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n646_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n827_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n647_), .B1(new_n835_), .B2(new_n830_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n826_), .A2(new_n834_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n634_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n588_), .A2(new_n840_), .A3(new_n509_), .A4(new_n637_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n637_), .A2(new_n509_), .A3(new_n579_), .A4(new_n587_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT113), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n843_), .A3(KEYINPUT54), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(KEYINPUT113), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n282_), .B1(new_n839_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n653_), .A2(new_n371_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n332_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT59), .B1(new_n849_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n847_), .B1(new_n838_), .B2(new_n634_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n282_), .A4(new_n851_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n795_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n833_), .B(new_n647_), .C1(new_n835_), .C2(new_n830_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n688_), .B1(new_n860_), .B2(new_n826_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n283_), .B(new_n852_), .C1(new_n861_), .C2(new_n847_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n855_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n849_), .A2(KEYINPUT59), .A3(new_n852_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(KEYINPUT118), .A3(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n857_), .A2(new_n700_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G113gat), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n509_), .A2(G113gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n862_), .B2(new_n868_), .ZN(G1340gat));
  AOI21_X1  g668(.A(new_n588_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n588_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(KEYINPUT60), .B2(new_n871_), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n870_), .A2(new_n871_), .B1(new_n862_), .B2(new_n873_), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n857_), .A2(new_n688_), .A3(new_n865_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G127gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n849_), .A2(new_n230_), .A3(new_n688_), .A4(new_n852_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(KEYINPUT119), .A3(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1342gat));
  OAI21_X1  g681(.A(new_n228_), .B1(new_n862_), .B2(new_n646_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT120), .Z(new_n884_));
  NAND4_X1  g683(.A1(new_n857_), .A2(new_n865_), .A3(G134gat), .A4(new_n696_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1343gat));
  NAND4_X1  g685(.A1(new_n849_), .A2(new_n371_), .A3(new_n333_), .A4(new_n714_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n509_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT121), .B(G141gat), .Z(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n588_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n219_), .ZN(G1345gat));
  NOR2_X1   g691(.A1(new_n887_), .A2(new_n634_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT61), .B(G155gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  INV_X1    g694(.A(G162gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n887_), .B2(new_n646_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT122), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n887_), .A2(new_n896_), .A3(new_n695_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1347gat));
  NAND3_X1  g699(.A1(new_n334_), .A2(new_n653_), .A3(new_n372_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n854_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n700_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n903_), .B(G169gat), .C1(KEYINPUT123), .C2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(KEYINPUT123), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT22), .B(G169gat), .Z(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n903_), .B2(new_n908_), .ZN(G1348gat));
  NAND2_X1  g708(.A1(new_n902_), .A2(new_n589_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n302_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT124), .B(G176gat), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n910_), .B2(new_n913_), .ZN(G1349gat));
  NAND2_X1  g713(.A1(new_n902_), .A2(new_n688_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n317_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT125), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n902_), .A2(KEYINPUT126), .A3(new_n688_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n915_), .B2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n918_), .B2(new_n920_), .ZN(G1350gat));
  NAND4_X1  g720(.A1(new_n902_), .A2(new_n393_), .A3(new_n395_), .A4(new_n647_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n854_), .A2(new_n695_), .A3(new_n901_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n394_), .ZN(G1351gat));
  NOR4_X1   g723(.A1(new_n854_), .A2(new_n443_), .A3(new_n332_), .A4(new_n714_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n700_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(KEYINPUT127), .B2(new_n352_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT127), .B(G197gat), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n589_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n350_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n346_), .B2(new_n930_), .ZN(G1353gat));
  NAND2_X1  g731(.A1(new_n925_), .A2(new_n688_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n936_), .B1(new_n933_), .B2(new_n934_), .ZN(G1354gat));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n925_), .A2(new_n938_), .A3(new_n647_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n925_), .A2(new_n696_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n938_), .ZN(G1355gat));
endmodule


