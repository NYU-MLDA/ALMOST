//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT4), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G113gat), .B(G120gat), .Z(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT77), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n210_), .B1(new_n214_), .B2(KEYINPUT77), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT84), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n223_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT83), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n228_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT83), .ZN(new_n231_));
  OR2_X1    g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT3), .ZN(new_n233_));
  AND4_X1   g032(.A1(new_n225_), .A2(new_n229_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT82), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(new_n236_), .B2(new_n232_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT3), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT81), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT82), .B(new_n238_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n220_), .B1(new_n234_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n232_), .A2(KEYINPUT79), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n238_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n248_), .A3(new_n226_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n219_), .B(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n218_), .B2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n206_), .B(new_n215_), .C1(new_n245_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT97), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n252_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n225_), .A2(new_n229_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n237_), .B2(new_n243_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n258_), .B2(new_n220_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n259_), .A2(KEYINPUT97), .A3(new_n206_), .A4(new_n215_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n215_), .B1(new_n245_), .B2(new_n252_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n214_), .B(new_n256_), .C1(new_n258_), .C2(new_n220_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT4), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G225gat), .A2(G233gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT96), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT98), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT98), .A4(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n205_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n271_), .A2(new_n272_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n205_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n255_), .A2(new_n260_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT89), .B(G204gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(G197gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(KEYINPUT21), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n283_), .B2(KEYINPUT21), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288_));
  INV_X1    g087(.A(G197gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT88), .B1(new_n289_), .B2(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT88), .ZN(new_n291_));
  INV_X1    g090(.A(G204gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(G197gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n282_), .A2(new_n289_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n288_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n285_), .B1(new_n287_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT90), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(G197gat), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT21), .B1(new_n303_), .B2(new_n294_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n304_), .B(new_n286_), .C1(KEYINPUT21), .C2(new_n283_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT90), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n285_), .ZN(new_n307_));
  OR2_X1    g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(KEYINPUT24), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT75), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n308_), .A2(KEYINPUT24), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT25), .B(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320_));
  INV_X1    g119(.A(G190gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT26), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G190gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n319_), .B(new_n322_), .C1(new_n323_), .C2(new_n320_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n311_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G176gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(G169gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G169gat), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n326_), .B(new_n329_), .C1(new_n330_), .C2(new_n327_), .ZN(new_n331_));
  OR2_X1    g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n314_), .A2(new_n332_), .A3(new_n315_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n309_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n299_), .A2(new_n307_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT20), .ZN(new_n338_));
  INV_X1    g137(.A(new_n302_), .ZN(new_n339_));
  OAI21_X1  g138(.A(G197gat), .B1(new_n339_), .B2(new_n300_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(G197gat), .B2(G204gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n284_), .A2(KEYINPUT21), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n284_), .B1(new_n341_), .B2(new_n288_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(new_n304_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n333_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n314_), .A2(new_n332_), .A3(KEYINPUT94), .A4(new_n315_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n330_), .A2(new_n326_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(new_n309_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n323_), .A2(new_n319_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n351_), .A2(new_n316_), .A3(new_n317_), .A4(new_n310_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n338_), .B1(new_n345_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT19), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n336_), .A2(new_n337_), .A3(new_n354_), .A4(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n336_), .A2(new_n357_), .A3(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT95), .ZN(new_n360_));
  INV_X1    g159(.A(new_n335_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n298_), .A2(KEYINPUT90), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n306_), .B1(new_n305_), .B2(new_n285_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n353_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n338_), .B1(new_n365_), .B2(new_n298_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n357_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n358_), .B1(new_n360_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n336_), .A2(new_n356_), .A3(new_n354_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n345_), .B2(new_n353_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n299_), .A2(new_n307_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n361_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n379_), .B2(new_n356_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(new_n374_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n280_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n262_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(new_n205_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n264_), .A2(new_n265_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n261_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT99), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n384_), .B(KEYINPUT99), .C1(new_n261_), .C2(new_n385_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n279_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n275_), .A2(KEYINPUT33), .A3(new_n276_), .A4(new_n278_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n368_), .A2(new_n373_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n372_), .B(new_n358_), .C1(new_n360_), .C2(new_n367_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n382_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT93), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT29), .B1(new_n245_), .B2(new_n252_), .ZN(new_n400_));
  INV_X1    g199(.A(G228gat), .ZN(new_n401_));
  INV_X1    g200(.A(G233gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n405_), .A2(new_n378_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n345_), .B1(new_n259_), .B2(KEYINPUT29), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n400_), .A2(new_n298_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(KEYINPUT91), .A3(new_n403_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n406_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n399_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT85), .B(KEYINPUT87), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G22gat), .B(G50gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n245_), .A2(new_n252_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NOR4_X1   g223(.A1(new_n245_), .A2(new_n252_), .A3(KEYINPUT29), .A4(new_n420_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n417_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n420_), .B1(new_n259_), .B2(KEYINPUT29), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n422_), .A2(new_n423_), .A3(new_n421_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n416_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n413_), .B(KEYINPUT92), .Z(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n412_), .B2(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n405_), .A2(new_n378_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT91), .B1(new_n410_), .B2(new_n403_), .ZN(new_n434_));
  AOI211_X1 g233(.A(new_n407_), .B(new_n404_), .C1(new_n400_), .C2(new_n298_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT93), .A3(new_n413_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n415_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n412_), .A2(new_n431_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n433_), .B(new_n431_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n430_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n398_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n372_), .B(new_n376_), .C1(new_n379_), .C2(new_n356_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT27), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT100), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n395_), .B2(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT95), .B(new_n359_), .C1(new_n379_), .C2(new_n357_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n372_), .B1(new_n449_), .B2(new_n358_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT100), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n452_));
  AOI22_X1  g251(.A1(new_n448_), .A2(new_n451_), .B1(new_n397_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n280_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n444_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(G15gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT30), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n459_), .B1(new_n325_), .B2(new_n334_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462_));
  INV_X1    g261(.A(G43gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n325_), .A2(new_n459_), .A3(new_n334_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n464_), .B1(new_n468_), .B2(new_n460_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n215_), .B(KEYINPUT31), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT78), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT31), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n215_), .B(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(KEYINPUT78), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n467_), .B(new_n469_), .C1(new_n472_), .C2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n469_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n396_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n452_), .B1(new_n482_), .B2(new_n450_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n446_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n450_), .B2(KEYINPUT100), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n395_), .A2(new_n447_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n483_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n274_), .A2(new_n279_), .A3(new_n480_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n442_), .A3(new_n438_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT102), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT102), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n453_), .A2(new_n443_), .A3(new_n491_), .A4(new_n488_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n456_), .A2(new_n481_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT34), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT35), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G85gat), .ZN(new_n499_));
  INV_X1    g298(.A(G92gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  INV_X1    g306(.A(G99gat), .ZN(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n503_), .B1(new_n506_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT8), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n515_), .B(new_n503_), .C1(new_n506_), .C2(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT10), .B(G99gat), .Z(new_n518_));
  AOI21_X1  g317(.A(new_n506_), .B1(new_n509_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT65), .B(G92gat), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT66), .B(new_n520_), .C1(new_n521_), .C2(new_n499_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n502_), .B1(new_n501_), .B2(KEYINPUT9), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n500_), .A2(KEYINPUT65), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n500_), .A2(KEYINPUT65), .ZN(new_n526_));
  OAI21_X1  g325(.A(G85gat), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT66), .B1(new_n527_), .B2(new_n520_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n519_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n517_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G43gat), .B(G50gat), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n498_), .B1(new_n530_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n535_), .B(KEYINPUT15), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n530_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n496_), .A2(KEYINPUT35), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n538_), .B(new_n540_), .C1(KEYINPUT70), .C2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(KEYINPUT70), .B(new_n498_), .C1(new_n530_), .C2(new_n536_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n540_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n543_), .B(new_n544_), .C1(new_n545_), .C2(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(KEYINPUT71), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(KEYINPUT36), .B2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(KEYINPUT36), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n542_), .A2(new_n546_), .A3(KEYINPUT71), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n550_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n494_), .B1(new_n554_), .B2(new_n560_), .ZN(new_n561_));
  AOI211_X1 g360(.A(KEYINPUT37), .B(new_n559_), .C1(new_n551_), .C2(new_n553_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT73), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G183gat), .B(G211gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572_));
  INV_X1    g371(.A(G1gat), .ZN(new_n573_));
  INV_X1    g372(.A(G8gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT14), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G1gat), .B(G8gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(KEYINPUT67), .ZN(new_n581_));
  INV_X1    g380(.A(G57gat), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(G64gat), .ZN(new_n583_));
  INV_X1    g382(.A(G64gat), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(G57gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n581_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT11), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(G57gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(G64gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT67), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n587_), .A3(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G71gat), .B(G78gat), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n590_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(KEYINPUT11), .ZN(new_n596_));
  AOI211_X1 g395(.A(KEYINPUT68), .B(new_n587_), .C1(new_n586_), .C2(new_n590_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT67), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT67), .B1(new_n588_), .B2(new_n589_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT11), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT68), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n594_), .A3(KEYINPUT11), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n580_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n571_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n570_), .B2(new_n569_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n563_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT64), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n596_), .A2(new_n597_), .A3(new_n593_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n602_), .A2(new_n603_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n530_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n598_), .A2(new_n604_), .A3(new_n529_), .A4(new_n517_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(KEYINPUT12), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n605_), .A2(new_n620_), .A3(new_n530_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n614_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n617_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n618_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n614_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(G120gat), .B(G148gat), .Z(new_n627_));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n623_), .A2(new_n626_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT13), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n631_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n536_), .A2(new_n578_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n539_), .A2(new_n578_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n536_), .B(new_n578_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n641_), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n642_), .A2(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(G113gat), .B(G141gat), .Z(new_n647_));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n646_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n639_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n493_), .A2(new_n611_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n280_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n655_), .A2(G1gat), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n658_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT38), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n559_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n493_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n610_), .A3(new_n652_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G1gat), .B1(new_n667_), .B2(new_n656_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n659_), .A2(KEYINPUT38), .A3(new_n660_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n663_), .A2(new_n668_), .A3(new_n669_), .ZN(G1324gat));
  NAND3_X1  g469(.A1(new_n654_), .A2(new_n574_), .A3(new_n487_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT104), .Z(new_n672_));
  OAI21_X1  g471(.A(G8gat), .B1(new_n667_), .B2(new_n453_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n674_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n672_), .A2(KEYINPUT40), .A3(new_n675_), .A4(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1325gat));
  OAI21_X1  g480(.A(G15gat), .B1(new_n667_), .B2(new_n481_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT41), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n655_), .A2(G15gat), .A3(new_n481_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1326gat));
  OR3_X1    g484(.A1(new_n655_), .A2(G22gat), .A3(new_n443_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n667_), .A2(new_n443_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n688_));
  AND3_X1   g487(.A1(new_n687_), .A2(G22gat), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n687_), .B2(G22gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(G1327gat));
  NOR2_X1   g490(.A1(new_n664_), .A2(new_n610_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n492_), .A2(new_n490_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n480_), .B1(new_n444_), .B2(new_n455_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n652_), .B(new_n692_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT106), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n438_), .A2(new_n442_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n656_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n487_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n482_), .A2(new_n450_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n700_), .A2(new_n393_), .A3(new_n390_), .A4(new_n392_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n701_), .B2(new_n382_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n481_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n492_), .A2(new_n490_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n652_), .A4(new_n692_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n696_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n280_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n493_), .B2(new_n563_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n664_), .B(new_n494_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n705_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n610_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n652_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT44), .B1(new_n714_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n719_), .B(new_n716_), .C1(new_n710_), .C2(new_n713_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n280_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n709_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  XNOR2_X1  g522(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n453_), .A2(G36gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n696_), .A2(new_n707_), .A3(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n728_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n696_), .A2(new_n707_), .A3(new_n730_), .A4(new_n726_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n711_), .B1(new_n705_), .B2(new_n712_), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT43), .B(new_n563_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n717_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n719_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n714_), .A2(KEYINPUT44), .A3(new_n717_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n487_), .A3(new_n737_), .ZN(new_n738_));
  AOI211_X1 g537(.A(new_n725_), .B(new_n732_), .C1(G36gat), .C2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(G36gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n732_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n724_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1329gat));
  XOR2_X1   g542(.A(KEYINPUT109), .B(G43gat), .Z(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n708_), .B2(new_n480_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n481_), .A2(new_n463_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n721_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(G1330gat));
  INV_X1    g548(.A(G50gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n721_), .B2(new_n697_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n697_), .A2(new_n750_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT110), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n708_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT111), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n718_), .A2(new_n720_), .A3(new_n443_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n757_), .B(new_n754_), .C1(new_n758_), .C2(new_n750_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1331gat));
  NAND4_X1  g559(.A1(new_n666_), .A2(new_n610_), .A3(new_n651_), .A4(new_n639_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n656_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n639_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n611_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT112), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n493_), .A2(new_n650_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n280_), .A2(new_n582_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n767_), .B2(new_n768_), .ZN(G1332gat));
  OAI21_X1  g568(.A(G64gat), .B1(new_n761_), .B2(new_n453_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT48), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n487_), .A2(new_n584_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n767_), .B2(new_n772_), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n761_), .B2(new_n481_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT49), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n481_), .A2(G71gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n767_), .B2(new_n776_), .ZN(G1334gat));
  OAI21_X1  g576(.A(G78gat), .B1(new_n761_), .B2(new_n443_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT50), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n443_), .A2(G78gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT113), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n767_), .B2(new_n781_), .ZN(G1335gat));
  AND3_X1   g581(.A1(new_n766_), .A2(new_n639_), .A3(new_n692_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n499_), .A3(new_n280_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n639_), .A2(new_n651_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(new_n610_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n714_), .A2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n280_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n788_), .B2(new_n499_), .ZN(G1336gat));
  AOI21_X1  g588(.A(G92gat), .B1(new_n783_), .B2(new_n487_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n453_), .A2(new_n521_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n787_), .B2(new_n791_), .ZN(G1337gat));
  NAND2_X1  g591(.A1(new_n480_), .A2(new_n518_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT114), .B1(new_n783_), .B2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n787_), .A2(new_n480_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n508_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n795_), .B(new_n798_), .C1(new_n796_), .C2(new_n508_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n783_), .A2(new_n509_), .A3(new_n697_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n714_), .A2(new_n697_), .A3(new_n786_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(G106gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n804_), .B2(G106gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT53), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n803_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n637_), .A2(new_n651_), .A3(new_n638_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT116), .B(new_n813_), .C1(new_n611_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n815_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n817_), .A2(new_n610_), .A3(new_n563_), .A4(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n814_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n631_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n619_), .A2(new_n614_), .A3(new_n621_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n622_), .B1(KEYINPUT55), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n824_), .B(new_n614_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT56), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n828_), .B(new_n821_), .C1(new_n823_), .C2(new_n825_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n827_), .A2(new_n650_), .A3(new_n632_), .A4(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n646_), .A2(new_n649_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n649_), .B1(new_n644_), .B2(new_n641_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n643_), .A2(new_n640_), .A3(new_n645_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n665_), .B1(new_n830_), .B2(new_n837_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n838_), .A2(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(KEYINPUT57), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n827_), .A2(new_n632_), .A3(new_n836_), .A4(new_n829_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n712_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n841_), .A2(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n843_), .B2(new_n712_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n839_), .B(new_n840_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n820_), .B1(new_n849_), .B2(new_n715_), .ZN(new_n850_));
  NOR4_X1   g649(.A1(new_n487_), .A2(new_n697_), .A3(new_n481_), .A4(new_n656_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853_), .B2(new_n650_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n843_), .A2(new_n712_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT117), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n846_), .A3(new_n845_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n838_), .B(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n610_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT59), .B(new_n851_), .C1(new_n862_), .C2(new_n820_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n856_), .A2(KEYINPUT118), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT118), .B1(new_n856_), .B2(new_n863_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n650_), .A2(G113gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n854_), .B1(new_n866_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n763_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n853_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n763_), .B1(new_n856_), .B2(new_n863_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n869_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n853_), .B2(new_n610_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n610_), .A2(new_n875_), .A3(G127gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n875_), .B2(G127gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n874_), .B1(new_n866_), .B2(new_n877_), .ZN(G1342gat));
  AOI21_X1  g677(.A(G134gat), .B1(new_n853_), .B2(new_n665_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n712_), .A2(G134gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n866_), .B2(new_n880_), .ZN(G1343gat));
  NOR4_X1   g680(.A1(new_n487_), .A2(new_n443_), .A3(new_n656_), .A4(new_n480_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT120), .B1(new_n850_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n885_), .B(new_n882_), .C1(new_n862_), .C2(new_n820_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n651_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT121), .B(G141gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1344gat));
  AOI21_X1  g688(.A(new_n763_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n890_));
  INV_X1    g689(.A(G148gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1345gat));
  AOI21_X1  g691(.A(new_n715_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n893_), .B(new_n895_), .ZN(G1346gat));
  NAND2_X1  g695(.A1(new_n884_), .A2(new_n886_), .ZN(new_n897_));
  INV_X1    g696(.A(G162gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n665_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n563_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1347gat));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n453_), .A2(new_n489_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n650_), .B(new_n903_), .C1(new_n862_), .C2(new_n820_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G169gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n905_), .B2(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(KEYINPUT62), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n904_), .A2(KEYINPUT122), .A3(new_n908_), .A4(G169gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n906_), .A2(new_n907_), .A3(new_n909_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n850_), .A2(new_n453_), .A3(new_n489_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n912_), .B(new_n903_), .C1(new_n862_), .C2(new_n820_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n330_), .B(new_n650_), .C1(new_n913_), .C2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n910_), .A2(new_n916_), .ZN(G1348gat));
  OAI21_X1  g716(.A(new_n639_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919_));
  INV_X1    g718(.A(new_n850_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n903_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n763_), .A2(new_n326_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n919_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n911_), .A2(KEYINPUT124), .A3(new_n922_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n918_), .A2(new_n326_), .B1(new_n924_), .B2(new_n925_), .ZN(G1349gat));
  AOI21_X1  g725(.A(G183gat), .B1(new_n911_), .B2(new_n610_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n921_), .A2(KEYINPUT123), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n914_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n715_), .A2(new_n319_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n927_), .B1(new_n929_), .B2(new_n930_), .ZN(G1350gat));
  NAND2_X1  g730(.A1(new_n665_), .A2(new_n323_), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n932_), .B(KEYINPUT125), .Z(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n563_), .B1(new_n928_), .B2(new_n914_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n321_), .ZN(G1351gat));
  NOR3_X1   g735(.A1(new_n698_), .A2(new_n453_), .A3(new_n480_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n920_), .A2(new_n650_), .A3(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g738(.A1(new_n920_), .A2(new_n639_), .A3(new_n937_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n282_), .B1(KEYINPUT126), .B2(new_n292_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n940_), .B2(new_n943_), .ZN(G1353gat));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n715_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n920_), .A2(new_n945_), .A3(new_n937_), .A4(new_n946_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n937_), .B(new_n946_), .C1(new_n862_), .C2(new_n820_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(KEYINPUT127), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1354gat));
  INV_X1    g751(.A(G218gat), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n920_), .A2(new_n953_), .A3(new_n665_), .A4(new_n937_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n920_), .A2(new_n712_), .A3(new_n937_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n954_), .B1(new_n956_), .B2(new_n953_), .ZN(G1355gat));
endmodule


