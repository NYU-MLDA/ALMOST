//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_,
    new_n588_, new_n590_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  AND3_X1   g004(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  AOI211_X1 g007(.A(new_n204_), .B(new_n206_), .C1(new_n207_), .C2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  MUX2_X1   g011(.A(new_n212_), .B(new_n210_), .S(KEYINPUT23), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(new_n212_), .B2(KEYINPUT23), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT22), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n221_), .A2(KEYINPUT81), .A3(G169gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT81), .B1(new_n221_), .B2(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n223_), .B(new_n224_), .C1(KEYINPUT22), .C2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n220_), .B(new_n205_), .C1(new_n222_), .C2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n214_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G71gat), .B(G99gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT82), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT31), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n241_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G155gat), .A2(G162gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G141gat), .A2(G148gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT3), .Z(new_n250_));
  NAND2_X1  g049(.A1(G141gat), .A2(G148gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT2), .Z(new_n252_));
  OAI211_X1 g051(.A(new_n246_), .B(new_n248_), .C1(new_n250_), .C2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n247_), .B1(KEYINPUT1), .B2(new_n246_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(KEYINPUT1), .B2(new_n246_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n249_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT29), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G228gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(G78gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G106gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n261_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(G211gat), .B(G218gat), .Z(new_n268_));
  INV_X1    g067(.A(KEYINPUT21), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G197gat), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(G204gat), .ZN(new_n272_));
  AOI211_X1 g071(.A(new_n269_), .B(new_n268_), .C1(KEYINPUT84), .C2(new_n272_), .ZN(new_n273_));
  MUX2_X1   g072(.A(new_n270_), .B(new_n267_), .S(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275_));
  INV_X1    g074(.A(new_n258_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G22gat), .B(G50gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n266_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n266_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT18), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n209_), .A2(new_n216_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n213_), .A2(new_n290_), .A3(new_n219_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G169gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n224_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n205_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n290_), .B1(new_n213_), .B2(new_n219_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n289_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n274_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n300_), .B1(new_n299_), .B2(new_n274_), .ZN(new_n302_));
  OAI221_X1 g101(.A(KEYINPUT20), .B1(new_n274_), .B2(new_n228_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT88), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT19), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n274_), .A2(new_n228_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(KEYINPUT20), .C1(new_n274_), .C2(new_n299_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n304_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n288_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n303_), .A2(new_n306_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT88), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n315_), .A2(new_n287_), .A3(new_n307_), .A4(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n276_), .A2(new_n235_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n234_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n233_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n258_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(KEYINPUT90), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT4), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n319_), .A2(new_n326_), .A3(new_n258_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n325_), .B(new_n327_), .C1(new_n321_), .C2(new_n326_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n324_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT89), .B(KEYINPUT0), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n331_), .A2(KEYINPUT91), .A3(KEYINPUT33), .A4(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n324_), .A2(new_n328_), .A3(new_n336_), .A4(new_n330_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT33), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n323_), .B(new_n327_), .C1(new_n321_), .C2(new_n326_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(KEYINPUT92), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(KEYINPUT92), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT33), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n337_), .A2(new_n341_), .B1(new_n346_), .B2(new_n339_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n313_), .A2(new_n316_), .A3(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n331_), .A2(new_n336_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT94), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n339_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n331_), .A2(KEYINPUT94), .A3(new_n336_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n309_), .A2(new_n306_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(KEYINPUT32), .A3(new_n287_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n307_), .A2(new_n310_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n287_), .A2(KEYINPUT32), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n315_), .A3(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n348_), .A2(KEYINPUT93), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT93), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n313_), .A2(new_n316_), .A3(new_n362_), .A4(new_n347_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n283_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n287_), .B1(new_n358_), .B2(new_n315_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n311_), .A2(new_n288_), .A3(new_n312_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n353_), .A2(new_n282_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n355_), .A2(new_n288_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n316_), .A2(KEYINPUT27), .A3(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n369_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n245_), .B1(new_n364_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n369_), .A2(new_n282_), .A3(new_n372_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT96), .ZN(new_n376_));
  INV_X1    g175(.A(new_n353_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT96), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n369_), .A2(new_n378_), .A3(new_n282_), .A4(new_n372_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n244_), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G29gat), .B(G36gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G43gat), .B(G50gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT15), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G15gat), .B(G22gat), .ZN(new_n386_));
  INV_X1    g185(.A(G1gat), .ZN(new_n387_));
  INV_X1    g186(.A(G8gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT14), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G1gat), .B(G8gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n385_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n384_), .B(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G229gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n395_), .B(new_n392_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G113gat), .B(G141gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(G169gat), .B(G197gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n404_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT97), .B1(new_n381_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT97), .ZN(new_n409_));
  INV_X1    g208(.A(new_n407_), .ZN(new_n410_));
  AOI211_X1 g209(.A(new_n409_), .B(new_n410_), .C1(new_n374_), .C2(new_n380_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G230gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G64gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G57gat), .ZN(new_n415_));
  INV_X1    g214(.A(G57gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G64gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT68), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT11), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n416_), .A2(G64gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n414_), .A2(G57gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT68), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT11), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G78gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n421_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT69), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT11), .B(new_n428_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT10), .B(G99gat), .Z(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G85gat), .B(G92gat), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT9), .ZN(new_n440_));
  INV_X1    g239(.A(G85gat), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  OR3_X1    g241(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT9), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT6), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n438_), .A2(new_n440_), .A3(new_n443_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT7), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT64), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT65), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT65), .A4(new_n455_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT66), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT67), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n448_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n445_), .A2(new_n447_), .A3(new_n463_), .A4(new_n465_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n439_), .B1(new_n461_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT8), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n458_), .A2(new_n448_), .A3(new_n459_), .A4(new_n460_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n439_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT8), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n450_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n435_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n435_), .B2(new_n476_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n471_), .A2(new_n475_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n430_), .A2(new_n432_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT69), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n481_), .A2(new_n449_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n413_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n449_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n487_), .A2(KEYINPUT12), .A3(new_n432_), .A4(new_n430_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n413_), .B1(new_n435_), .B2(new_n476_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n470_), .A2(KEYINPUT8), .B1(new_n472_), .B2(new_n474_), .ZN(new_n490_));
  OAI22_X1  g289(.A1(new_n490_), .A2(new_n450_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT71), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT12), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n488_), .B(new_n489_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n486_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G120gat), .B(G148gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT5), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G176gat), .B(G204gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n486_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT13), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n502_), .B(new_n504_), .C1(KEYINPUT72), .C2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n408_), .A2(new_n411_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT34), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n487_), .A2(new_n385_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n516_), .B1(new_n517_), .B2(KEYINPUT73), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n476_), .A2(new_n384_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n517_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n522_), .B2(new_n518_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G190gat), .B(G218gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT36), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(KEYINPUT74), .Z(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(KEYINPUT37), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n523_), .A2(KEYINPUT75), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT75), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n520_), .B(new_n537_), .C1(new_n518_), .C2(new_n522_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT76), .B1(new_n539_), .B2(new_n527_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT76), .ZN(new_n541_));
  AOI211_X1 g340(.A(new_n541_), .B(new_n528_), .C1(new_n536_), .C2(new_n538_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n533_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n535_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G127gat), .B(G155gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT16), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G183gat), .B(G211gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT77), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n392_), .B(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n552_), .B1(new_n555_), .B2(new_n482_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n482_), .B2(new_n555_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT78), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n550_), .A2(new_n551_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n435_), .ZN(new_n561_));
  AOI211_X1 g360(.A(new_n552_), .B(new_n560_), .C1(new_n555_), .C2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n555_), .B2(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n546_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n513_), .A2(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n566_), .A2(G1gat), .A3(new_n377_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n543_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n571_), .A2(new_n564_), .A3(new_n512_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n381_), .A2(new_n407_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(G1gat), .B1(new_n574_), .B2(new_n377_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n570_), .A3(new_n575_), .ZN(G1324gat));
  NAND2_X1  g375(.A1(new_n369_), .A2(new_n372_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n388_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT39), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n577_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(G8gat), .ZN(new_n581_));
  AOI211_X1 g380(.A(KEYINPUT39), .B(new_n388_), .C1(new_n573_), .C2(new_n577_), .ZN(new_n582_));
  OAI22_X1  g381(.A1(new_n566_), .A2(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(G1325gat));
  AOI21_X1  g384(.A(new_n238_), .B1(new_n573_), .B2(new_n244_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT41), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n244_), .A2(new_n238_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n587_), .B1(new_n566_), .B2(new_n588_), .ZN(G1326gat));
  INV_X1    g388(.A(G22gat), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n573_), .B2(new_n283_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT42), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n283_), .A2(new_n590_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n566_), .B2(new_n593_), .ZN(G1327gat));
  INV_X1    g393(.A(new_n564_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n512_), .A2(new_n595_), .A3(new_n410_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT43), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n381_), .B2(new_n546_), .ZN(new_n598_));
  AOI211_X1 g397(.A(KEYINPUT43), .B(new_n545_), .C1(new_n374_), .C2(new_n380_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT44), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT44), .B(new_n596_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n353_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(G29gat), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n543_), .A2(new_n595_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n513_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(G29gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n353_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT100), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n609_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1328gat));
  NAND3_X1  g413(.A1(new_n602_), .A2(new_n577_), .A3(new_n603_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G36gat), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n408_), .A2(new_n512_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n411_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n577_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(G36gat), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n606_), .A4(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT45), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT45), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n513_), .A2(new_n623_), .A3(new_n606_), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n616_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT46), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n616_), .A2(KEYINPUT46), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1329gat));
  NAND4_X1  g429(.A1(new_n602_), .A2(G43gat), .A3(new_n244_), .A4(new_n603_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n617_), .A2(new_n244_), .A3(new_n618_), .A4(new_n606_), .ZN(new_n632_));
  INV_X1    g431(.A(G43gat), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n632_), .A2(KEYINPUT101), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT101), .B1(new_n632_), .B2(new_n633_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT47), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT47), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(new_n631_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1330gat));
  NAND3_X1  g439(.A1(new_n602_), .A2(new_n283_), .A3(new_n603_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G50gat), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n282_), .A2(G50gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT102), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n607_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(G1331gat));
  AOI211_X1 g445(.A(new_n407_), .B(new_n511_), .C1(new_n374_), .C2(new_n380_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(new_n595_), .A3(new_n543_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT103), .B(G57gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n353_), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT104), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n647_), .A2(new_n565_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G57gat), .B1(new_n652_), .B2(new_n353_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1332gat));
  AOI21_X1  g453(.A(new_n414_), .B1(new_n648_), .B2(new_n577_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT48), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n414_), .A3(new_n577_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1333gat));
  INV_X1    g457(.A(G71gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n648_), .B2(new_n244_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT49), .Z(new_n661_));
  NAND3_X1  g460(.A1(new_n652_), .A2(new_n659_), .A3(new_n244_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1334gat));
  AOI21_X1  g462(.A(new_n263_), .B1(new_n648_), .B2(new_n283_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT50), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n652_), .A2(new_n263_), .A3(new_n283_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1335gat));
  NAND2_X1  g466(.A1(new_n647_), .A2(new_n606_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n441_), .B1(new_n668_), .B2(new_n377_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n669_), .A2(new_n670_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n598_), .A2(new_n599_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n511_), .A2(new_n595_), .A3(new_n407_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n377_), .A2(new_n441_), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n671_), .B(new_n672_), .C1(new_n675_), .C2(new_n676_), .ZN(G1336gat));
  OAI21_X1  g476(.A(new_n442_), .B1(new_n668_), .B2(new_n619_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n678_), .A2(new_n679_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n619_), .A2(new_n442_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n680_), .B(new_n681_), .C1(new_n675_), .C2(new_n682_), .ZN(G1337gat));
  NAND3_X1  g482(.A1(new_n673_), .A2(new_n244_), .A3(new_n674_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G99gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n668_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n436_), .A3(new_n244_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT107), .B(KEYINPUT51), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(G1338gat));
  NAND3_X1  g489(.A1(new_n686_), .A2(new_n437_), .A3(new_n283_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n283_), .B(new_n674_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT52), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G106gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G106gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g496(.A(new_n404_), .B1(new_n400_), .B2(new_n397_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n397_), .B2(new_n396_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n505_), .A2(new_n406_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n407_), .A2(new_n504_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT56), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT55), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n496_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT71), .B1(new_n485_), .B2(KEYINPUT12), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n707_), .A2(KEYINPUT55), .A3(new_n488_), .A4(new_n489_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n478_), .A2(new_n479_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n707_), .A2(new_n710_), .A3(new_n711_), .A4(new_n488_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n711_), .A3(new_n488_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n412_), .B1(new_n713_), .B2(KEYINPUT109), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n709_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n702_), .B1(new_n715_), .B2(new_n503_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n488_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT109), .B1(new_n717_), .B2(new_n480_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n413_), .A3(new_n712_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n704_), .A3(new_n708_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(KEYINPUT56), .A3(new_n501_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n701_), .B1(new_n716_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n700_), .B1(new_n722_), .B2(KEYINPUT110), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n724_), .B(new_n701_), .C1(new_n716_), .C2(new_n721_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n543_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT57), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n721_), .A2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n720_), .A2(KEYINPUT111), .A3(KEYINPUT56), .A4(new_n501_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n716_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n504_), .A2(new_n406_), .A3(new_n699_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT58), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(KEYINPUT58), .A3(new_n733_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n546_), .A3(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT57), .B(new_n543_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n728_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n564_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n595_), .A2(new_n410_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n511_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT108), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n511_), .A2(new_n747_), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n742_), .B1(new_n749_), .B2(new_n545_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n747_), .B1(new_n511_), .B2(new_n744_), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT108), .B(new_n743_), .C1(new_n508_), .C2(new_n510_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n545_), .B(new_n742_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n750_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n741_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n376_), .A2(new_n244_), .A3(new_n379_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n353_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(KEYINPUT113), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT113), .B(KEYINPUT59), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n377_), .B1(new_n741_), .B2(new_n756_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n759_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n763_), .A2(new_n410_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(G113gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n760_), .A2(KEYINPUT112), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n765_), .A2(new_n770_), .A3(new_n759_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n407_), .A2(new_n768_), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n767_), .A2(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(G1340gat));
  NOR3_X1   g573(.A1(new_n763_), .A2(new_n511_), .A3(new_n766_), .ZN(new_n775_));
  INV_X1    g574(.A(G120gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n511_), .B2(KEYINPUT60), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(KEYINPUT60), .B2(new_n776_), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n775_), .A2(new_n776_), .B1(new_n772_), .B2(new_n778_), .ZN(G1341gat));
  INV_X1    g578(.A(G127gat), .ZN(new_n780_));
  NOR4_X1   g579(.A1(new_n763_), .A2(new_n766_), .A3(new_n780_), .A4(new_n564_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n770_), .B1(new_n765_), .B2(new_n759_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n755_), .B1(new_n740_), .B2(new_n564_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n784_), .A2(KEYINPUT112), .A3(new_n377_), .A4(new_n758_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n783_), .A2(new_n785_), .A3(new_n564_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n786_), .B2(G127gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n769_), .A2(new_n595_), .A3(new_n771_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(KEYINPUT114), .A3(new_n780_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n781_), .B1(new_n787_), .B2(new_n789_), .ZN(G1342gat));
  INV_X1    g589(.A(G134gat), .ZN(new_n791_));
  NOR4_X1   g590(.A1(new_n763_), .A2(new_n766_), .A3(new_n791_), .A4(new_n545_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n783_), .A2(new_n785_), .A3(new_n543_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G134gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n769_), .A2(new_n571_), .A3(new_n771_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT115), .A3(new_n791_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n792_), .B1(new_n795_), .B2(new_n797_), .ZN(G1343gat));
  NAND2_X1  g597(.A1(new_n757_), .A2(new_n353_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n619_), .A2(new_n283_), .A3(new_n245_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n407_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT116), .B(G141gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1344gat));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n512_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT117), .B(G148gat), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n805_), .B(new_n806_), .Z(G1345gat));
  NAND2_X1  g606(.A1(new_n801_), .A2(new_n595_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT61), .B(G155gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  NOR2_X1   g609(.A1(new_n543_), .A2(G162gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n801_), .A2(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n799_), .A2(new_n545_), .A3(new_n800_), .ZN(new_n813_));
  INV_X1    g612(.A(G162gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n812_), .B(KEYINPUT118), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1347gat));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n784_), .A2(new_n619_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n245_), .A2(new_n283_), .A3(new_n353_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n822_), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n784_), .A2(KEYINPUT121), .A3(new_n619_), .A4(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n407_), .A2(new_n292_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT122), .Z(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n821_), .A2(new_n822_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT119), .B1(new_n832_), .B2(new_n410_), .ZN(new_n833_));
  NOR4_X1   g632(.A1(new_n784_), .A2(new_n410_), .A3(new_n619_), .A4(new_n825_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n225_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n833_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n831_), .B1(new_n839_), .B2(new_n840_), .ZN(G1348gat));
  NAND3_X1  g640(.A1(new_n828_), .A2(new_n224_), .A3(new_n512_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G176gat), .B1(new_n832_), .B2(new_n511_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1349gat));
  NOR2_X1   g643(.A1(new_n564_), .A2(new_n207_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(new_n845_), .C1(new_n823_), .C2(new_n826_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n217_), .B1(new_n832_), .B2(new_n564_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(G1350gat));
  NAND3_X1  g650(.A1(new_n828_), .A2(new_n571_), .A3(new_n208_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n545_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n218_), .ZN(G1351gat));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855_));
  AND4_X1   g654(.A1(new_n370_), .A2(new_n757_), .A3(new_n577_), .A4(new_n245_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n407_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(new_n271_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n856_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n407_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n271_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(G1352gat));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G204gat), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT125), .B(G204gat), .Z(new_n864_));
  NAND2_X1  g663(.A1(new_n856_), .A2(new_n512_), .ZN(new_n865_));
  MUX2_X1   g664(.A(new_n863_), .B(new_n864_), .S(new_n865_), .Z(G1353gat));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n867_));
  INV_X1    g666(.A(G211gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n595_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT126), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n868_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n856_), .A2(new_n870_), .B1(KEYINPUT127), .B2(new_n871_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n871_), .A2(KEYINPUT127), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1354gat));
  INV_X1    g673(.A(G218gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n856_), .A2(new_n875_), .A3(new_n571_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n856_), .A2(new_n546_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n875_), .ZN(G1355gat));
endmodule


