//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT67), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n202_), .A2(new_n203_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OR3_X1    g009(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT7), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(KEYINPUT7), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G85gat), .B(G92gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n217_), .B2(KEYINPUT66), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n219_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n223_), .A2(new_n214_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT10), .B(G99gat), .ZN(new_n226_));
  OAI221_X1 g025(.A(new_n224_), .B1(KEYINPUT9), .B2(new_n225_), .C1(G106gat), .C2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n210_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT12), .ZN(new_n230_));
  INV_X1    g029(.A(new_n228_), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n231_), .A2(new_n210_), .A3(KEYINPUT12), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G230gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT64), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(new_n236_), .B2(new_n229_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G120gat), .B(G148gat), .ZN(new_n239_));
  INV_X1    g038(.A(G204gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT5), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G176gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n238_), .B(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT13), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(KEYINPUT13), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(KEYINPUT68), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G1gat), .A2(G8gat), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n250_), .A2(KEYINPUT14), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT75), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G15gat), .B(G22gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G1gat), .B(G8gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G231gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(new_n210_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G127gat), .B(G155gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G183gat), .B(G211gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT17), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(KEYINPUT17), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n260_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(KEYINPUT77), .Z(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n266_), .B2(new_n260_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G190gat), .B(G218gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G134gat), .ZN(new_n273_));
  INV_X1    g072(.A(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT36), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n275_), .A2(new_n276_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT69), .B(G43gat), .ZN(new_n280_));
  INV_X1    g079(.A(G50gat), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n280_), .A2(new_n281_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT70), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT15), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n228_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G232gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT34), .Z(new_n294_));
  INV_X1    g093(.A(KEYINPUT35), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n228_), .A2(new_n287_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(KEYINPUT71), .A3(new_n228_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n292_), .A2(new_n296_), .A3(new_n297_), .A4(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n294_), .A2(new_n295_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT73), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n299_), .A2(KEYINPUT74), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT74), .B1(new_n299_), .B2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n292_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n300_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT72), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n277_), .B(new_n279_), .C1(new_n306_), .C2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n309_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n311_), .A2(new_n276_), .A3(new_n275_), .A4(new_n305_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT37), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT37), .B1(new_n310_), .B2(new_n312_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n249_), .A2(new_n271_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT91), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G211gat), .A2(G218gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT91), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT21), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(G204gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n240_), .A2(G197gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n327_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n240_), .A2(G197gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(G204gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT90), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .A4(KEYINPUT21), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT90), .B1(new_n329_), .B2(G204gat), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n340_), .A2(KEYINPUT21), .B1(new_n335_), .B2(new_n336_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n327_), .B(KEYINPUT92), .C1(new_n339_), .C2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n337_), .B1(G197gat), .B2(new_n240_), .ZN(new_n344_));
  OAI22_X1  g143(.A1(new_n344_), .A2(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n338_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT92), .B1(new_n346_), .B2(new_n327_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n334_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G169gat), .ZN(new_n351_));
  INV_X1    g150(.A(G176gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT24), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358_));
  INV_X1    g157(.A(G190gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(KEYINPUT26), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT25), .B(G183gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G190gat), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n360_), .B(new_n361_), .C1(new_n362_), .C2(new_n358_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n355_), .A2(new_n354_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n357_), .A2(new_n363_), .A3(new_n368_), .A4(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G169gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n353_), .B1(new_n371_), .B2(new_n352_), .ZN(new_n372_));
  OR2_X1    g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n366_), .A2(new_n373_), .A3(new_n367_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n327_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT92), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n342_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(KEYINPUT93), .A3(new_n334_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n350_), .A2(new_n377_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n333_), .B1(new_n380_), .B2(new_n342_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n387_));
  AND4_X1   g186(.A1(new_n386_), .A2(new_n369_), .A3(new_n367_), .A4(new_n366_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n356_), .B1(new_n362_), .B2(new_n361_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n374_), .B(KEYINPUT96), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n389_), .A2(new_n390_), .B1(new_n391_), .B2(new_n372_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n384_), .B1(new_n385_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n387_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n388_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n372_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n348_), .A2(new_n398_), .A3(KEYINPUT97), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n383_), .A2(KEYINPUT20), .A3(new_n393_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(KEYINPUT94), .Z(new_n402_));
  XOR2_X1   g201(.A(new_n402_), .B(KEYINPUT19), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT18), .B(G64gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G92gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT93), .B1(new_n381_), .B2(new_n334_), .ZN(new_n409_));
  AOI211_X1 g208(.A(new_n349_), .B(new_n333_), .C1(new_n380_), .C2(new_n342_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n376_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n403_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n385_), .A2(new_n392_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(KEYINPUT20), .A3(new_n412_), .A4(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n404_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(KEYINPUT20), .A3(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n403_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n393_), .A2(new_n399_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n418_), .A2(KEYINPUT20), .A3(new_n412_), .A4(new_n383_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n408_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n415_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n408_), .B1(new_n404_), .B2(new_n414_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n415_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n425_), .A2(KEYINPUT106), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(KEYINPUT106), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT2), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n431_));
  OAI22_X1  g230(.A1(new_n429_), .A2(new_n430_), .B1(new_n431_), .B2(KEYINPUT87), .ZN(new_n432_));
  INV_X1    g231(.A(G141gat), .ZN(new_n433_));
  INV_X1    g232(.A(G148gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n433_), .B(new_n434_), .C1(new_n435_), .C2(KEYINPUT3), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n431_), .B(KEYINPUT87), .C1(G141gat), .C2(G148gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n432_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT88), .B(KEYINPUT2), .ZN(new_n439_));
  INV_X1    g238(.A(new_n429_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT89), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n430_), .A2(KEYINPUT88), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n430_), .A2(KEYINPUT88), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n442_), .B(new_n429_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n438_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n433_), .A2(new_n434_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(new_n429_), .C1(new_n451_), .C2(new_n448_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT86), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n448_), .A2(new_n451_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(new_n440_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n454_), .A4(new_n452_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n450_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(KEYINPUT29), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT28), .ZN(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(KEYINPUT29), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n468_), .B(new_n469_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n348_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(G228gat), .A3(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G22gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G78gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n470_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n467_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n466_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n376_), .B(KEYINPUT30), .Z(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G227gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n485_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT84), .B(G113gat), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G120gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(G127gat), .B(G134gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT84), .B(G113gat), .ZN(new_n493_));
  INV_X1    g292(.A(G120gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n491_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G99gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n489_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G1gat), .B(G29gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G57gat), .B(G85gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  OR2_X1    g305(.A1(new_n496_), .A2(new_n497_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT98), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n507_), .B(new_n508_), .C1(new_n462_), .C2(new_n509_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n446_), .A2(new_n449_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n498_), .B1(new_n511_), .B2(KEYINPUT98), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT98), .B1(new_n511_), .B2(KEYINPUT99), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n510_), .B(KEYINPUT4), .C1(new_n512_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G225gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT100), .B(KEYINPUT4), .Z(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n462_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n510_), .B(new_n515_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n506_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n506_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n501_), .A2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n428_), .A2(new_n482_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n415_), .A2(new_n423_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n510_), .B1(new_n513_), .B2(new_n512_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT102), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n510_), .B(KEYINPUT102), .C1(new_n512_), .C2(new_n513_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n516_), .A3(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n514_), .A2(new_n518_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n534_), .B(KEYINPUT33), .C1(new_n516_), .C2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n506_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n519_), .A2(new_n520_), .A3(new_n506_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT33), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n519_), .A2(new_n520_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT33), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n529_), .A2(new_n538_), .A3(new_n540_), .A4(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n417_), .A2(new_n419_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n404_), .B2(new_n414_), .ZN(new_n546_));
  OAI22_X1  g345(.A1(new_n545_), .A2(new_n546_), .B1(new_n521_), .B2(new_n539_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT103), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n524_), .B(KEYINPUT103), .C1(new_n546_), .C2(new_n545_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n543_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n481_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT104), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n425_), .A2(new_n524_), .A3(new_n481_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(KEYINPUT104), .A3(new_n481_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n501_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n558_), .A2(KEYINPUT105), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT105), .B1(new_n558_), .B2(new_n559_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n528_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n287_), .B(KEYINPUT79), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n257_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT80), .ZN(new_n565_));
  INV_X1    g364(.A(new_n257_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n289_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n563_), .A2(new_n257_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n351_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n329_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT81), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n573_), .B(new_n577_), .Z(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT82), .Z(new_n579_));
  AND2_X1   g378(.A1(new_n562_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n319_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n317_), .A2(new_n318_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n583_), .A2(G1gat), .A3(new_n525_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT107), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT38), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT107), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n584_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n310_), .A2(new_n312_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT108), .Z(new_n592_));
  INV_X1    g391(.A(new_n247_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n578_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n592_), .A2(new_n595_), .A3(new_n271_), .A4(new_n562_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n525_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n590_), .A3(new_n597_), .ZN(G1324gat));
  INV_X1    g397(.A(new_n428_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n583_), .A2(G8gat), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT109), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  OAI221_X1 g401(.A(G8gat), .B1(new_n601_), .B2(new_n602_), .C1(new_n596_), .C2(new_n599_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(KEYINPUT109), .A2(KEYINPUT39), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g406(.A(G15gat), .B1(new_n596_), .B2(new_n559_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT41), .Z(new_n609_));
  OR2_X1    g408(.A1(new_n559_), .A2(G15gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n583_), .B2(new_n610_), .ZN(G1326gat));
  OAI21_X1  g410(.A(G22gat), .B1(new_n596_), .B2(new_n481_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT110), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT42), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n581_), .A2(new_n482_), .A3(new_n582_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n614_), .B1(G22gat), .B2(new_n615_), .ZN(G1327gat));
  NOR2_X1   g415(.A1(new_n592_), .A2(new_n271_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n580_), .A3(new_n247_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT113), .ZN(new_n619_));
  AOI21_X1  g418(.A(G29gat), .B1(new_n619_), .B2(new_n524_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT111), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n551_), .A2(KEYINPUT104), .A3(new_n481_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT104), .B1(new_n551_), .B2(new_n481_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n555_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n622_), .B1(new_n625_), .B2(new_n501_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n558_), .A2(KEYINPUT105), .A3(new_n559_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n527_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT43), .B1(new_n628_), .B2(new_n316_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  INV_X1    g429(.A(new_n315_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n313_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n562_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n595_), .A2(new_n270_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n621_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  AOI211_X1 g436(.A(KEYINPUT111), .B(new_n635_), .C1(new_n629_), .C2(new_n633_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT112), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT112), .ZN(new_n642_));
  NOR4_X1   g441(.A1(new_n637_), .A2(new_n638_), .A3(new_n642_), .A4(KEYINPUT44), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n634_), .A2(new_n636_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n640_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n644_), .A2(new_n525_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n620_), .B1(new_n647_), .B2(G29gat), .ZN(G1328gat));
  NOR2_X1   g447(.A1(KEYINPUT115), .A2(KEYINPUT46), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT115), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n646_), .A2(new_n599_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT114), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT114), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n653_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(G36gat), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n619_), .A2(new_n659_), .A3(new_n428_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT45), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n649_), .B(new_n652_), .C1(new_n658_), .C2(new_n661_), .ZN(new_n662_));
  AND4_X1   g461(.A1(new_n650_), .A2(new_n658_), .A3(new_n651_), .A4(new_n661_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  NOR2_X1   g463(.A1(new_n644_), .A2(new_n646_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(G43gat), .A3(new_n501_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n619_), .A2(new_n501_), .ZN(new_n667_));
  INV_X1    g466(.A(G43gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g470(.A(G50gat), .B1(new_n619_), .B2(new_n482_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n481_), .A2(new_n281_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n665_), .B2(new_n673_), .ZN(G1331gat));
  NOR2_X1   g473(.A1(new_n249_), .A2(new_n628_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n579_), .A2(new_n270_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n592_), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G57gat), .B1(new_n677_), .B2(new_n525_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n247_), .A2(new_n578_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n562_), .A2(new_n271_), .A3(new_n316_), .A4(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n680_), .A2(G57gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n525_), .B2(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT116), .Z(G1332gat));
  OAI21_X1  g482(.A(G64gat), .B1(new_n677_), .B2(new_n599_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT48), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n599_), .A2(G64gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n680_), .B2(new_n686_), .ZN(G1333gat));
  OAI21_X1  g486(.A(G71gat), .B1(new_n677_), .B2(new_n559_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT49), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n559_), .A2(G71gat), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT117), .Z(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n680_), .B2(new_n691_), .ZN(G1334gat));
  OAI21_X1  g491(.A(G78gat), .B1(new_n677_), .B2(new_n481_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT50), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n680_), .A2(G78gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n481_), .B2(new_n695_), .ZN(G1335gat));
  AND3_X1   g495(.A1(new_n675_), .A2(new_n594_), .A3(new_n617_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n524_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n679_), .A2(new_n270_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT118), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n634_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n524_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n698_), .B1(G85gat), .B2(new_n702_), .ZN(G1336gat));
  AOI21_X1  g502(.A(G92gat), .B1(new_n697_), .B2(new_n428_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT119), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n701_), .A2(G92gat), .A3(new_n428_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1337gat));
  NAND2_X1  g506(.A1(new_n701_), .A2(new_n501_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n559_), .A2(new_n226_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n708_), .A2(G99gat), .B1(new_n697_), .B2(new_n709_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g510(.A(new_n465_), .B1(new_n701_), .B2(new_n482_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT52), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n697_), .A2(new_n465_), .A3(new_n482_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g515(.A1(new_n676_), .A2(new_n316_), .A3(new_n247_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(KEYINPUT120), .B2(KEYINPUT54), .ZN(new_n718_));
  NAND2_X1  g517(.A1(KEYINPUT120), .A2(KEYINPUT54), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT121), .Z(new_n720_));
  XNOR2_X1  g519(.A(new_n718_), .B(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n237_), .B(KEYINPUT55), .Z(new_n722_));
  NOR2_X1   g521(.A1(new_n233_), .A2(new_n236_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n243_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT56), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n238_), .A2(new_n243_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n578_), .A3(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n568_), .A2(new_n569_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n730_));
  MUX2_X1   g529(.A(new_n573_), .B(new_n730_), .S(new_n576_), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n244_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n592_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT57), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n592_), .A2(new_n733_), .A3(KEYINPUT57), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n726_), .A2(new_n727_), .A3(new_n731_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT58), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n632_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n721_), .B1(new_n741_), .B2(new_n271_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n599_), .A2(new_n524_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n559_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(new_n481_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G113gat), .B1(new_n746_), .B2(new_n578_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT59), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n742_), .A2(KEYINPUT59), .A3(new_n481_), .A4(new_n744_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  XOR2_X1   g550(.A(KEYINPUT122), .B(G113gat), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n579_), .A2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT123), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n747_), .B1(new_n751_), .B2(new_n754_), .ZN(G1340gat));
  XOR2_X1   g554(.A(KEYINPUT124), .B(G120gat), .Z(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n247_), .B2(KEYINPUT60), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n746_), .B(new_n758_), .C1(KEYINPUT60), .C2(new_n757_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n249_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n757_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT125), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT125), .B(new_n759_), .C1(new_n760_), .C2(new_n757_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1341gat));
  AOI21_X1  g564(.A(G127gat), .B1(new_n746_), .B2(new_n271_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n270_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g567(.A(new_n592_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G134gat), .B1(new_n746_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n632_), .A2(G134gat), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT126), .Z(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n751_), .B2(new_n772_), .ZN(G1343gat));
  AND2_X1   g572(.A1(new_n742_), .A2(new_n559_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n743_), .A2(new_n481_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n594_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(new_n433_), .ZN(G1344gat));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n249_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(new_n434_), .ZN(G1345gat));
  NOR2_X1   g579(.A1(new_n776_), .A2(new_n270_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT61), .B(G155gat), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT127), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n781_), .B(new_n783_), .ZN(G1346gat));
  NOR3_X1   g583(.A1(new_n776_), .A2(new_n274_), .A3(new_n316_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n774_), .A2(new_n769_), .A3(new_n775_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n274_), .B2(new_n786_), .ZN(G1347gat));
  AND2_X1   g586(.A1(new_n742_), .A2(new_n481_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n526_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(new_n428_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n578_), .A3(new_n371_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n788_), .A2(new_n578_), .A3(new_n789_), .A4(new_n428_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(G169gat), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT62), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n792_), .A2(new_n794_), .A3(new_n797_), .ZN(G1348gat));
  NAND3_X1  g597(.A1(new_n791_), .A2(new_n352_), .A3(new_n593_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n790_), .A2(new_n428_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G176gat), .B1(new_n800_), .B2(new_n249_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1349gat));
  NAND3_X1  g601(.A1(new_n791_), .A2(new_n271_), .A3(new_n361_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G183gat), .B1(new_n800_), .B2(new_n270_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1350gat));
  NAND3_X1  g604(.A1(new_n791_), .A2(new_n769_), .A3(new_n362_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G190gat), .B1(new_n800_), .B2(new_n316_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1351gat));
  NOR3_X1   g607(.A1(new_n599_), .A2(new_n524_), .A3(new_n481_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n774_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n594_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(new_n329_), .ZN(G1352gat));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n249_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(new_n240_), .ZN(G1353gat));
  NOR2_X1   g613(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n815_));
  AND2_X1   g614(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n816_));
  NOR4_X1   g615(.A1(new_n810_), .A2(new_n270_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n774_), .A2(new_n809_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n271_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n819_), .B2(new_n815_), .ZN(G1354gat));
  AOI21_X1  g619(.A(G218gat), .B1(new_n818_), .B2(new_n769_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n810_), .A2(new_n316_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(G218gat), .B2(new_n822_), .ZN(G1355gat));
endmodule


