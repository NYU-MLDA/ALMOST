//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n977_, new_n978_, new_n979_, new_n980_, new_n982_,
    new_n983_;
  XOR2_X1   g000(.A(G197gat), .B(G204gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G228gat), .A2(G233gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(KEYINPUT93), .Z(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT88), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n222_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT89), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n217_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n220_), .A2(new_n221_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n214_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT90), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n214_), .A2(KEYINPUT90), .A3(new_n229_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT91), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n228_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n228_), .B(KEYINPUT92), .C1(new_n237_), .C2(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n227_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n211_), .B(new_n213_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G78gat), .B(G106gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT94), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n227_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n243_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT91), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n238_), .B(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(new_n236_), .A3(new_n232_), .A4(new_n235_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT92), .B1(new_n254_), .B2(new_n228_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n250_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n210_), .B1(new_n256_), .B2(KEYINPUT29), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n212_), .A2(KEYINPUT93), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n246_), .B(new_n249_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n244_), .A2(new_n260_), .A3(new_n245_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G22gat), .B(G50gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n244_), .A2(new_n245_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT28), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n268_), .B2(new_n261_), .ZN(new_n269_));
  OAI211_X1 g068(.A(KEYINPUT95), .B(new_n259_), .C1(new_n266_), .C2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n246_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n248_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT95), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n265_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(new_n271_), .A3(new_n248_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT96), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n271_), .B(new_n280_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n275_), .A2(new_n247_), .A3(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(G15gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT30), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT25), .B(G183gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT81), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(G169gat), .B2(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n296_), .A2(new_n298_), .A3(KEYINPUT24), .A4(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(G183gat), .B2(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n303_), .B1(new_n308_), .B2(new_n302_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n296_), .A2(new_n298_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n301_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n302_), .A2(G183gat), .A3(G190gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT84), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n306_), .A2(KEYINPUT23), .A3(new_n307_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n315_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT22), .B(G169gat), .Z(new_n320_));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n294_), .A2(KEYINPUT22), .ZN(new_n323_));
  AOI21_X1  g122(.A(G176gat), .B1(new_n323_), .B2(KEYINPUT83), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n299_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n314_), .B1(new_n319_), .B2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G71gat), .B(G99gat), .Z(new_n328_));
  XOR2_X1   g127(.A(KEYINPUT85), .B(G43gat), .Z(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NOR2_X1   g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n322_), .A2(new_n324_), .B1(G169gat), .B2(G176gat), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n317_), .A2(new_n318_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n315_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(new_n314_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n290_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n327_), .A2(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n314_), .A3(new_n332_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n289_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT31), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n285_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n337_), .A2(new_n340_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n349_), .A2(KEYINPUT86), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n353_));
  AOI211_X1 g152(.A(KEYINPUT87), .B(new_n347_), .C1(new_n337_), .C2(new_n340_), .ZN(new_n354_));
  OAI22_X1  g153(.A1(new_n348_), .A2(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n346_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n256_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT99), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n346_), .B(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(new_n250_), .C1(new_n255_), .C2(new_n251_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n365_), .A3(KEYINPUT4), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n256_), .A2(new_n369_), .A3(new_n361_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n366_), .A2(KEYINPUT100), .A3(new_n368_), .A4(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n368_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT100), .B1(new_n375_), .B2(new_n366_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n360_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT100), .ZN(new_n378_));
  INV_X1    g177(.A(new_n366_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n374_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n360_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n372_), .A4(new_n371_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n355_), .A2(new_n377_), .A3(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT19), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n317_), .A2(new_n318_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n313_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT97), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n317_), .A2(new_n318_), .B1(new_n312_), .B2(new_n311_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT97), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n396_), .A3(new_n301_), .ZN(new_n397_));
  OAI221_X1 g196(.A(new_n299_), .B1(G176gat), .B2(new_n320_), .C1(new_n309_), .C2(new_n315_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n210_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT20), .B1(new_n327_), .B2(new_n211_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n390_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n301_), .B1(new_n395_), .B2(KEYINPUT97), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n391_), .A2(KEYINPUT97), .A3(new_n313_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n210_), .B(new_n398_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n211_), .A2(new_n327_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n390_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT20), .A4(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n388_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n401_), .A2(new_n388_), .A3(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  INV_X1    g211(.A(new_n388_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n404_), .A2(KEYINPUT20), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n414_), .A2(KEYINPUT102), .B1(new_n211_), .B2(new_n327_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT102), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n404_), .A2(new_n416_), .A3(KEYINPUT20), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n406_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n399_), .A2(new_n400_), .A3(new_n390_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n413_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n410_), .A2(KEYINPUT27), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n411_), .A2(new_n412_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n284_), .A2(new_n383_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT104), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT104), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n284_), .A2(new_n383_), .A3(new_n425_), .A4(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n414_), .A2(KEYINPUT102), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n405_), .A3(new_n417_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n419_), .B1(new_n428_), .B2(new_n390_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n388_), .A2(KEYINPUT32), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT103), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT103), .ZN(new_n432_));
  INV_X1    g231(.A(new_n430_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n432_), .B(new_n433_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n377_), .A2(new_n382_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n401_), .A2(new_n407_), .A3(new_n430_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n362_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n360_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n370_), .A2(new_n367_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n366_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n411_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n382_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n373_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(KEYINPUT33), .A3(new_n381_), .A4(new_n380_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n438_), .A2(new_n448_), .A3(new_n284_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n420_), .A2(new_n421_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n410_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n412_), .B1(new_n451_), .B2(new_n408_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n450_), .A2(new_n382_), .A3(new_n377_), .A4(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n273_), .A2(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n355_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n424_), .A2(new_n426_), .B1(new_n449_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT65), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT64), .ZN(new_n458_));
  NAND2_X1  g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT64), .A3(new_n459_), .ZN(new_n464_));
  AOI21_X1  g263(.A(G106gat), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G85gat), .ZN(new_n466_));
  INV_X1    g265(.A(G92gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G85gat), .A2(G92gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT9), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G99gat), .A3(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n470_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n457_), .B1(new_n465_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n460_), .A2(new_n461_), .A3(new_n458_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT64), .B1(new_n463_), .B2(new_n459_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n470_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n483_), .A3(KEYINPUT65), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n487_));
  INV_X1    g286(.A(G99gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n479_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n473_), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n486_), .B(new_n489_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n493_));
  AND2_X1   g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n468_), .A2(KEYINPUT66), .A3(new_n469_), .ZN(new_n497_));
  AND4_X1   g296(.A1(new_n485_), .A2(new_n492_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n496_), .A2(new_n497_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n485_), .B1(new_n499_), .B2(new_n492_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n478_), .B(new_n484_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT67), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G29gat), .B(G36gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G43gat), .B(G50gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n492_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n496_), .A2(new_n497_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT8), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n499_), .A2(new_n485_), .A3(new_n492_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT67), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n478_), .A4(new_n484_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n502_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT70), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n502_), .A2(new_n516_), .A3(KEYINPUT70), .A4(new_n509_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT68), .B(KEYINPUT15), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n506_), .A2(new_n508_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n501_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT34), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT35), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n521_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(KEYINPUT35), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(KEYINPUT69), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n501_), .A2(new_n535_), .A3(new_n525_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n532_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G190gat), .B(G218gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT71), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT36), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n543_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n532_), .B(new_n549_), .C1(new_n533_), .C2(new_n538_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(KEYINPUT37), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(KEYINPUT73), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n554_));
  INV_X1    g353(.A(new_n537_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n533_), .B1(new_n521_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n530_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n554_), .B(new_n546_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(new_n550_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n502_), .A2(new_n516_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(KEYINPUT11), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(KEYINPUT11), .ZN(new_n571_));
  INV_X1    g370(.A(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n568_), .A2(KEYINPUT11), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n570_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n567_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n502_), .A2(new_n575_), .A3(new_n516_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n501_), .A2(KEYINPUT12), .A3(new_n576_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n580_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n583_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n566_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n587_), .A3(new_n566_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT13), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n590_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n588_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n575_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(G22gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n287_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G15gat), .A2(G22gat), .ZN(new_n601_));
  AND2_X1   g400(.A1(KEYINPUT74), .A2(G8gat), .ZN(new_n602_));
  NOR2_X1   g401(.A1(KEYINPUT74), .A2(G8gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  AOI221_X4 g403(.A(KEYINPUT75), .B1(new_n600_), .B2(new_n601_), .C1(new_n604_), .C2(KEYINPUT14), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(KEYINPUT14), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n601_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G1gat), .B(G8gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n605_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT14), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT74), .B(G8gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n614_), .B2(G1gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n608_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT75), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n607_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n610_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n598_), .B1(new_n612_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n575_), .B(new_n596_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n618_), .A3(new_n610_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n611_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT76), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n620_), .A2(new_n624_), .A3(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT16), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n628_), .A3(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT77), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n632_), .A2(new_n633_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n634_), .B(new_n637_), .C1(new_n624_), .C2(new_n620_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n636_), .A2(KEYINPUT78), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT78), .B1(new_n636_), .B2(new_n639_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n561_), .A2(new_n595_), .A3(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n509_), .B1(new_n612_), .B2(new_n619_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G229gat), .A2(G233gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n525_), .A2(new_n623_), .A3(new_n622_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT79), .ZN(new_n648_));
  INV_X1    g447(.A(new_n645_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n509_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n623_), .A2(new_n622_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n623_), .B2(new_n622_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT79), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n644_), .A2(new_n654_), .A3(new_n646_), .A4(new_n645_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G113gat), .B(G141gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G169gat), .B(G197gat), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n656_), .B(new_n657_), .Z(new_n658_));
  NAND4_X1  g457(.A1(new_n648_), .A2(new_n653_), .A3(new_n655_), .A4(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT80), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n653_), .A2(new_n655_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT80), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n648_), .A4(new_n658_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n648_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n658_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n456_), .A2(new_n643_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n436_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n671_), .A2(G1gat), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT38), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n559_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n456_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n595_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n636_), .A2(new_n639_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n669_), .A3(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n672_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n673_), .A2(new_n674_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n675_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1324gat));
  OR3_X1    g486(.A1(new_n671_), .A2(new_n422_), .A3(new_n614_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n450_), .A2(new_n452_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n681_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G8gat), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(KEYINPUT39), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(KEYINPUT39), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n694_), .B(new_n696_), .ZN(G1325gat));
  AOI21_X1  g496(.A(new_n287_), .B1(new_n681_), .B2(new_n355_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT41), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n670_), .A2(new_n287_), .A3(new_n355_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1326gat));
  AOI21_X1  g500(.A(new_n599_), .B1(new_n681_), .B2(new_n454_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT42), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n670_), .A2(new_n599_), .A3(new_n454_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1327gat));
  NOR2_X1   g504(.A1(new_n456_), .A2(new_n669_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n640_), .A2(new_n641_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n676_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n678_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n710_), .A2(G29gat), .A3(new_n672_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n456_), .B2(new_n561_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n449_), .A2(new_n455_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n454_), .A2(new_n689_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n425_), .B1(new_n714_), .B2(new_n383_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n426_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n558_), .A2(new_n550_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n554_), .B1(new_n539_), .B2(new_n546_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n560_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n551_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n717_), .A2(new_n718_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n712_), .A2(new_n723_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n678_), .A2(new_n642_), .A3(new_n669_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(KEYINPUT44), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n724_), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n724_), .B2(new_n725_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n436_), .A3(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT108), .ZN(new_n734_));
  OAI21_X1  g533(.A(G29gat), .B1(new_n733_), .B2(KEYINPUT108), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n711_), .B1(new_n734_), .B2(new_n735_), .ZN(G1328gat));
  INV_X1    g535(.A(new_n710_), .ZN(new_n737_));
  INV_X1    g536(.A(G36gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n689_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT45), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n731_), .A2(new_n422_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n730_), .A2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(KEYINPUT46), .B(new_n740_), .C1(new_n742_), .C2(new_n738_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  INV_X1    g543(.A(new_n740_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n738_), .B1(new_n730_), .B2(new_n741_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n747_), .ZN(G1329gat));
  AOI21_X1  g547(.A(G43gat), .B1(new_n737_), .B2(new_n355_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n730_), .A2(new_n732_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n355_), .A2(G43gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT47), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n750_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1330gat));
  AOI21_X1  g556(.A(G50gat), .B1(new_n737_), .B2(new_n454_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n751_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n454_), .A2(G50gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n595_), .A2(new_n668_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR4_X1   g562(.A1(new_n456_), .A2(new_n763_), .A3(new_n707_), .A4(new_n676_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n672_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n456_), .A2(new_n668_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n707_), .A2(new_n722_), .A3(new_n595_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT109), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(KEYINPUT109), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n436_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n767_), .B1(new_n774_), .B2(new_n766_), .ZN(G1332gat));
  OAI21_X1  g574(.A(G64gat), .B1(new_n765_), .B2(new_n422_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT48), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n422_), .A2(G64gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n770_), .B2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n771_), .A2(new_n780_), .A3(new_n355_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n764_), .B2(new_n355_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n783_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n784_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n781_), .B1(new_n787_), .B2(new_n788_), .ZN(G1334gat));
  OAI21_X1  g588(.A(G78gat), .B1(new_n765_), .B2(new_n284_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT50), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n284_), .A2(G78gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n770_), .B2(new_n792_), .ZN(G1335gat));
  NAND2_X1  g592(.A1(new_n762_), .A2(new_n707_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n724_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n672_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n768_), .A2(new_n678_), .A3(new_n707_), .A4(new_n676_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n466_), .A3(new_n436_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n796_), .B2(new_n422_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n467_), .A3(new_n689_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1337gat));
  INV_X1    g603(.A(new_n355_), .ZN(new_n805_));
  OAI21_X1  g604(.A(G99gat), .B1(new_n796_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n355_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n798_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n799_), .A2(new_n479_), .A3(new_n454_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n284_), .B(new_n794_), .C1(new_n712_), .C2(new_n723_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n479_), .B1(new_n813_), .B2(KEYINPUT112), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n794_), .B1(new_n712_), .B2(new_n723_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n815_), .B2(new_n454_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n724_), .A2(KEYINPUT112), .A3(new_n454_), .A4(new_n795_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G106gat), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n820_), .A2(new_n816_), .A3(new_n811_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n810_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT53), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n810_), .C1(new_n818_), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1339gat));
  NOR4_X1   g625(.A1(new_n454_), .A2(new_n672_), .A3(new_n689_), .A4(new_n805_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n679_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n645_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n644_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n831_), .A2(new_n666_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n592_), .B2(new_n588_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n586_), .B2(KEYINPUT114), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n836_), .B2(new_n586_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n579_), .A2(new_n582_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT12), .B1(new_n567_), .B2(new_n576_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n580_), .A2(new_n581_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n837_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AND4_X1   g641(.A1(KEYINPUT56), .A2(new_n839_), .A3(new_n565_), .A4(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n575_), .B1(new_n502_), .B2(new_n516_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n580_), .B(new_n581_), .C1(new_n844_), .C2(KEYINPUT12), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n566_), .B1(new_n845_), .B2(new_n837_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n839_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n668_), .B(new_n590_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n558_), .A2(new_n550_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n835_), .A2(new_n848_), .B1(new_n849_), .B2(new_n553_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n829_), .B(new_n830_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n835_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n559_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT117), .B1(new_n854_), .B2(KEYINPUT115), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n850_), .B2(new_n829_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n590_), .B(new_n834_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n721_), .A2(new_n551_), .B1(new_n859_), .B2(new_n858_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(KEYINPUT116), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n858_), .A2(new_n859_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n561_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n828_), .B1(new_n857_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n643_), .B2(new_n668_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n707_), .A2(new_n722_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n669_), .A4(new_n595_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n827_), .B1(new_n867_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G113gat), .B1(new_n874_), .B2(new_n668_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n830_), .B1(new_n854_), .B2(KEYINPUT117), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n829_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n879_), .A2(new_n852_), .B1(new_n865_), .B2(new_n862_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n876_), .B1(new_n880_), .B2(new_n642_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n868_), .A2(new_n871_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n857_), .A2(new_n866_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(KEYINPUT120), .A3(new_n707_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n827_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n827_), .A2(new_n886_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n887_), .A2(new_n888_), .A3(KEYINPUT59), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT121), .B1(new_n885_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n642_), .B1(new_n857_), .B2(new_n866_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n882_), .B1(new_n892_), .B2(KEYINPUT120), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n880_), .A2(new_n876_), .A3(new_n642_), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT121), .B(new_n889_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT118), .B1(new_n873_), .B2(KEYINPUT59), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n873_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n891_), .A2(new_n895_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n668_), .A2(G113gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n875_), .B1(new_n899_), .B2(new_n900_), .ZN(G1340gat));
  INV_X1    g700(.A(new_n895_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n890_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n873_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n678_), .B1(new_n904_), .B2(new_n896_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G120gat), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n595_), .A2(KEYINPUT60), .ZN(new_n907_));
  MUX2_X1   g706(.A(new_n907_), .B(KEYINPUT60), .S(G120gat), .Z(new_n908_));
  NAND2_X1  g707(.A1(new_n874_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n909_), .ZN(G1341gat));
  AOI21_X1  g709(.A(G127gat), .B1(new_n874_), .B2(new_n642_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n828_), .A2(G127gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n899_), .B2(new_n912_), .ZN(G1342gat));
  AOI21_X1  g712(.A(G134gat), .B1(new_n874_), .B2(new_n676_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n722_), .A2(G134gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n899_), .B2(new_n915_), .ZN(G1343gat));
  OAI21_X1  g715(.A(new_n882_), .B1(new_n880_), .B2(new_n828_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n284_), .A2(new_n355_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n672_), .A2(new_n689_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n669_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT122), .B(G141gat), .Z(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1344gat));
  NOR2_X1   g722(.A1(new_n920_), .A2(new_n595_), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g724(.A1(new_n920_), .A2(new_n707_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT61), .B(G155gat), .Z(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n920_), .B2(new_n561_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n559_), .A2(G162gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n920_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n422_), .A2(new_n436_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n355_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n454_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n885_), .A2(new_n668_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(G169gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n938_), .A2(new_n320_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n939_), .A2(new_n940_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(G1348gat));
  NAND2_X1  g743(.A1(new_n917_), .A2(new_n284_), .ZN(new_n945_));
  OR4_X1    g744(.A1(new_n295_), .A2(new_n945_), .A3(new_n595_), .A4(new_n936_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n885_), .A2(new_n678_), .A3(new_n937_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(KEYINPUT125), .A3(new_n295_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  INV_X1    g749(.A(new_n948_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(G176gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n947_), .B1(new_n949_), .B2(new_n952_), .ZN(G1349gat));
  NOR2_X1   g752(.A1(new_n679_), .A2(new_n291_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n885_), .A2(new_n937_), .A3(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(G183gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n642_), .A2(new_n355_), .A3(new_n935_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n945_), .B2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n955_), .A2(new_n958_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(KEYINPUT126), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n885_), .A2(new_n722_), .A3(new_n937_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(G190gat), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n885_), .A2(new_n292_), .A3(new_n676_), .A4(new_n937_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n962_), .A2(KEYINPUT127), .A3(new_n963_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(G1351gat));
  AND2_X1   g767(.A1(new_n917_), .A2(new_n918_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n935_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n970_), .A2(new_n669_), .ZN(new_n971_));
  INV_X1    g770(.A(G197gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1352gat));
  NOR2_X1   g772(.A1(new_n970_), .A2(new_n595_), .ZN(new_n974_));
  INV_X1    g773(.A(G204gat), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n974_), .B(new_n975_), .ZN(G1353gat));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n977_), .B1(new_n970_), .B2(new_n679_), .ZN(new_n978_));
  XOR2_X1   g777(.A(KEYINPUT63), .B(G211gat), .Z(new_n979_));
  NAND4_X1  g778(.A1(new_n969_), .A2(new_n828_), .A3(new_n935_), .A4(new_n979_), .ZN(new_n980_));
  AND2_X1   g779(.A1(new_n978_), .A2(new_n980_), .ZN(G1354gat));
  OAI21_X1  g780(.A(G218gat), .B1(new_n970_), .B2(new_n561_), .ZN(new_n982_));
  OR2_X1    g781(.A1(new_n559_), .A2(G218gat), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n982_), .B1(new_n970_), .B2(new_n983_), .ZN(G1355gat));
endmodule


