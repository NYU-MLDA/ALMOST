//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OR2_X1    g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G169gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT78), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n203_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n218_), .A2(KEYINPUT77), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(KEYINPUT77), .ZN(new_n220_));
  OAI21_X1  g019(.A(G190gat), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n218_), .A2(G190gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT76), .ZN(new_n223_));
  INV_X1    g022(.A(G183gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT25), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(G183gat), .A3(new_n227_), .ZN(new_n228_));
  AND4_X1   g027(.A1(new_n221_), .A2(new_n223_), .A3(new_n225_), .A4(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n208_), .B1(new_n217_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT80), .ZN(new_n232_));
  XOR2_X1   g031(.A(G71gat), .B(G99gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n230_), .B(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G127gat), .B(G134gat), .Z(new_n236_));
  XOR2_X1   g035(.A(G113gat), .B(G120gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n235_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G15gat), .B(G43gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT79), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n239_), .B(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT3), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G141gat), .A2(G148gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT2), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n250_), .B1(KEYINPUT1), .B2(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(KEYINPUT1), .B2(new_n252_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n245_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n256_), .A2(new_n247_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n249_), .A2(new_n253_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n238_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT88), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n258_), .B2(new_n238_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n249_), .A2(new_n253_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n255_), .A2(new_n257_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n238_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(new_n261_), .A3(new_n259_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n269_), .A3(KEYINPUT4), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G29gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G85gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT0), .B(G57gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n263_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n269_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n274_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n276_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n281_), .B1(new_n276_), .B2(new_n284_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n244_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G8gat), .B(G36gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT18), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G64gat), .B(G92gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT19), .ZN(new_n296_));
  XOR2_X1   g095(.A(G211gat), .B(G218gat), .Z(new_n297_));
  INV_X1    g096(.A(G197gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(G204gat), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT81), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(G204gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(KEYINPUT81), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n297_), .B1(new_n303_), .B2(KEYINPUT21), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT21), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT82), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n297_), .A2(KEYINPUT21), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(KEYINPUT83), .B2(new_n305_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n305_), .A2(KEYINPUT83), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n304_), .A2(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n313_), .B2(new_n230_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT25), .B(G183gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n214_), .A2(new_n216_), .A3(new_n315_), .A4(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n205_), .A2(KEYINPUT86), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n321_), .A3(new_n204_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n207_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(new_n312_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n296_), .B1(new_n314_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n312_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n313_), .A2(new_n230_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n296_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT20), .A4(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n294_), .B1(new_n327_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(new_n294_), .A3(new_n331_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(KEYINPUT87), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(KEYINPUT87), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n332_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n340_));
  INV_X1    g139(.A(new_n230_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(new_n312_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n342_), .B(new_n330_), .C1(new_n312_), .C2(new_n325_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT20), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n296_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT27), .B(new_n334_), .C1(new_n346_), .C2(new_n294_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n339_), .A2(new_n347_), .ZN(new_n348_));
  OR3_X1    g147(.A1(new_n266_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT28), .B1(new_n266_), .B2(KEYINPUT29), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G22gat), .B(G50gat), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n258_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n313_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(G228gat), .B(G233gat), .C1(new_n312_), .C2(new_n358_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G78gat), .B(G106gat), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n355_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT85), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n363_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT84), .A4(new_n362_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n372_), .B2(new_n355_), .ZN(new_n373_));
  AOI211_X1 g172(.A(KEYINPUT85), .B(new_n354_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n367_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n348_), .A2(new_n376_), .A3(KEYINPUT91), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n339_), .A2(new_n347_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n375_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n289_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n274_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n382_));
  AOI211_X1 g181(.A(new_n281_), .B(new_n382_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n285_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n286_), .A2(KEYINPUT33), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n337_), .A2(new_n332_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n337_), .A2(new_n332_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n385_), .B(new_n386_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n294_), .A2(KEYINPUT32), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n343_), .A2(new_n345_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n327_), .B2(new_n331_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT89), .B1(new_n288_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT89), .ZN(new_n395_));
  OAI221_X1 g194(.A(new_n395_), .B1(new_n391_), .B2(new_n392_), .C1(new_n286_), .C2(new_n287_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n389_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n376_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n348_), .A2(new_n399_), .A3(new_n288_), .A4(new_n375_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n375_), .A2(new_n339_), .A3(new_n347_), .A4(new_n288_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT90), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n244_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n381_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G29gat), .B(G36gat), .Z(new_n406_));
  XOR2_X1   g205(.A(G43gat), .B(G50gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G15gat), .B(G22gat), .ZN(new_n410_));
  INV_X1    g209(.A(G1gat), .ZN(new_n411_));
  INV_X1    g210(.A(G8gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT14), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G8gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n409_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G229gat), .A2(G233gat), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n408_), .B(KEYINPUT15), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n416_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n409_), .B(new_n416_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n418_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n419_), .A2(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G113gat), .B(G141gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(G169gat), .B(G197gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n424_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT12), .ZN(new_n430_));
  INV_X1    g229(.A(G85gat), .ZN(new_n431_));
  INV_X1    g230(.A(G92gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G85gat), .A2(G92gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT6), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(G99gat), .A3(G106gat), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441_));
  INV_X1    g240(.A(G99gat), .ZN(new_n442_));
  INV_X1    g241(.A(G106gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n435_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT67), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT8), .B1(new_n435_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n434_), .B1(new_n433_), .B2(KEYINPUT9), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n432_), .A2(KEYINPUT66), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT66), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G92gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n431_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n456_));
  OAI21_X1  g255(.A(new_n451_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT64), .B(G106gat), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n460_), .A2(new_n461_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  OAI221_X1 g262(.A(new_n435_), .B1(new_n448_), .B2(KEYINPUT8), .C1(new_n440_), .C2(new_n446_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n450_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G57gat), .B(G64gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G71gat), .B(G78gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT11), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n469_));
  INV_X1    g268(.A(new_n467_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n465_), .A2(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n449_), .A2(new_n447_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n473_), .A3(new_n464_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n430_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G230gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT12), .B1(new_n465_), .B2(new_n474_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n479_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G120gat), .B(G148gat), .Z(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G176gat), .B(G204gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n482_), .A2(new_n483_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n496_));
  NAND3_X1  g295(.A1(new_n490_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT70), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n500_), .A3(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n465_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n409_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n420_), .B2(new_n503_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G232gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT34), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT35), .Z(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(KEYINPUT71), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(KEYINPUT35), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n509_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT71), .B1(new_n505_), .B2(new_n508_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514_));
  XOR2_X1   g313(.A(G134gat), .B(G162gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(G190gat), .B(G218gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n514_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n517_), .A2(new_n514_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n519_), .B(new_n520_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n518_), .A2(KEYINPUT37), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT37), .B1(new_n518_), .B2(new_n521_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT73), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G127gat), .B(G155gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G183gat), .B(G211gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT17), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(KEYINPUT17), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n416_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n473_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n532_), .A2(new_n535_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT74), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n524_), .A2(new_n539_), .ZN(new_n540_));
  NOR4_X1   g339(.A1(new_n405_), .A2(new_n429_), .A3(new_n502_), .A4(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(KEYINPUT92), .Z(new_n542_));
  INV_X1    g341(.A(new_n288_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n411_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT38), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n518_), .A2(new_n521_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n405_), .A2(new_n548_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n502_), .A2(KEYINPUT93), .A3(new_n429_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT93), .B1(new_n502_), .B2(new_n429_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n550_), .A2(new_n538_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(G1gat), .B1(new_n553_), .B2(new_n288_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n544_), .A2(new_n545_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n546_), .A2(new_n554_), .A3(new_n555_), .ZN(G1324gat));
  NAND3_X1  g355(.A1(new_n542_), .A2(new_n412_), .A3(new_n379_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n553_), .A2(new_n348_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n559_), .B2(new_n412_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT94), .B(G8gat), .C1(new_n553_), .C2(new_n348_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(KEYINPUT39), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT39), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n558_), .B(new_n563_), .C1(new_n559_), .C2(new_n412_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n557_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT40), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n557_), .A2(new_n562_), .A3(KEYINPUT40), .A4(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(G1325gat));
  INV_X1    g368(.A(G15gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n542_), .A2(new_n570_), .A3(new_n244_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT97), .ZN(new_n572_));
  OAI21_X1  g371(.A(G15gat), .B1(new_n553_), .B2(new_n404_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT95), .B(KEYINPUT41), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n542_), .A2(new_n581_), .A3(new_n570_), .A4(new_n244_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n572_), .A2(new_n579_), .A3(new_n580_), .A4(new_n582_), .ZN(G1326gat));
  INV_X1    g382(.A(G22gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n375_), .B(KEYINPUT98), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n542_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G22gat), .B1(new_n553_), .B2(new_n585_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT42), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(KEYINPUT42), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n587_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT99), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n587_), .B(new_n593_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(G1327gat));
  NOR2_X1   g394(.A1(new_n405_), .A2(new_n429_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n502_), .A2(new_n539_), .A3(new_n547_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n598_), .A2(G29gat), .A3(new_n288_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT43), .B1(new_n405_), .B2(new_n524_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT43), .ZN(new_n601_));
  INV_X1    g400(.A(new_n524_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n376_), .A2(new_n397_), .B1(new_n401_), .B2(KEYINPUT90), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n244_), .B1(new_n603_), .B2(new_n400_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n601_), .B(new_n602_), .C1(new_n604_), .C2(new_n381_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n539_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n550_), .A2(new_n607_), .A3(new_n551_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT100), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(KEYINPUT44), .A3(new_n609_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n543_), .A3(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n614_), .A2(KEYINPUT101), .A3(G29gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT101), .B1(new_n614_), .B2(G29gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n599_), .B1(new_n615_), .B2(new_n616_), .ZN(G1328gat));
  XNOR2_X1  g416(.A(new_n379_), .B(KEYINPUT102), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(G36gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n598_), .A2(KEYINPUT45), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT45), .B1(new_n598_), .B2(new_n621_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n612_), .A2(new_n379_), .A3(new_n613_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(new_n620_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT46), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT46), .B(new_n624_), .C1(new_n625_), .C2(new_n620_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1329gat));
  NAND4_X1  g429(.A1(new_n612_), .A2(G43gat), .A3(new_n244_), .A4(new_n613_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n598_), .A2(new_n404_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(G43gat), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g433(.A1(new_n598_), .A2(G50gat), .A3(new_n585_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n612_), .A2(new_n375_), .A3(new_n613_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n636_), .B2(G50gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT103), .ZN(G1331gat));
  INV_X1    g437(.A(new_n502_), .ZN(new_n639_));
  NOR4_X1   g438(.A1(new_n405_), .A2(new_n428_), .A3(new_n639_), .A4(new_n540_), .ZN(new_n640_));
  INV_X1    g439(.A(G57gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n543_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n549_), .A2(new_n429_), .A3(new_n502_), .A4(new_n539_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(new_n543_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n647_), .B2(new_n641_), .ZN(G1332gat));
  INV_X1    g447(.A(G64gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n640_), .A2(new_n649_), .A3(new_n619_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n619_), .A3(new_n646_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT48), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n651_), .A2(new_n652_), .A3(G64gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n651_), .B2(G64gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n653_), .B2(new_n654_), .ZN(G1333gat));
  INV_X1    g454(.A(G71gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n640_), .A2(new_n656_), .A3(new_n244_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n244_), .A3(new_n646_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT49), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n658_), .A2(new_n659_), .A3(G71gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n658_), .B2(G71gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(G1334gat));
  INV_X1    g461(.A(G78gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n640_), .A2(new_n663_), .A3(new_n586_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n645_), .A2(new_n586_), .A3(new_n646_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n666_));
  AND3_X1   g465(.A1(new_n665_), .A2(G78gat), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n665_), .B2(G78gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(G1335gat));
  NOR2_X1   g468(.A1(new_n405_), .A2(new_n428_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n639_), .A2(new_n539_), .A3(new_n547_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n431_), .A3(new_n543_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n607_), .A2(new_n502_), .A3(new_n429_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(new_n543_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n677_), .B2(new_n431_), .ZN(G1336gat));
  AOI21_X1  g477(.A(G92gat), .B1(new_n673_), .B2(new_n379_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n618_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n676_), .B2(new_n680_), .ZN(G1337gat));
  NAND2_X1  g480(.A1(new_n244_), .A2(new_n460_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n672_), .A2(KEYINPUT106), .A3(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT106), .B1(new_n672_), .B2(new_n682_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n676_), .A2(new_n244_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n442_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT51), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n687_), .B(new_n689_), .Z(G1338gat));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n376_), .B(new_n675_), .C1(new_n600_), .C2(new_n605_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(new_n443_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n676_), .A2(new_n375_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(KEYINPUT110), .A3(G106gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n696_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n691_), .B(new_n698_), .C1(new_n692_), .C2(new_n443_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n375_), .A2(new_n670_), .A3(new_n461_), .A4(new_n671_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n699_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT53), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT53), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n697_), .A2(new_n705_), .A3(new_n699_), .A4(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1339gat));
  INV_X1    g506(.A(KEYINPUT54), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n539_), .A2(new_n429_), .A3(new_n498_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n539_), .A2(KEYINPUT111), .A3(new_n429_), .A4(new_n498_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n708_), .B1(new_n713_), .B2(new_n524_), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT54), .B(new_n602_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n421_), .A2(new_n417_), .A3(new_n423_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n427_), .B1(new_n422_), .B2(new_n418_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n424_), .A2(new_n427_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n492_), .A2(KEYINPUT115), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT115), .B1(new_n492_), .B2(new_n720_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n428_), .A2(new_n490_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT56), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n473_), .B1(new_n476_), .B2(new_n464_), .ZN(new_n726_));
  AND4_X1   g525(.A1(new_n473_), .A2(new_n450_), .A3(new_n464_), .A4(new_n463_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT12), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n481_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n728_), .A2(KEYINPUT55), .A3(new_n479_), .A4(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n480_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n479_), .A3(new_n729_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT113), .B(new_n732_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n489_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT112), .B1(new_n482_), .B2(KEYINPUT55), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT113), .B1(new_n742_), .B2(new_n732_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n725_), .B1(new_n739_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n732_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n747_), .A2(KEYINPUT56), .A3(new_n489_), .A4(new_n738_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n724_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n723_), .B1(new_n749_), .B2(KEYINPUT114), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n751_), .B(new_n724_), .C1(new_n744_), .C2(new_n748_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n547_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(KEYINPUT116), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT116), .B1(new_n753_), .B2(new_n754_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT57), .B(new_n547_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n490_), .A2(new_n720_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n524_), .B1(new_n759_), .B2(KEYINPUT58), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(KEYINPUT58), .B2(new_n759_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n761_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n755_), .A2(new_n756_), .A3(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n717_), .B1(new_n763_), .B2(new_n538_), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n404_), .B(new_n288_), .C1(new_n377_), .C2(new_n380_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT59), .ZN(new_n767_));
  INV_X1    g566(.A(new_n723_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n724_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n739_), .A2(new_n743_), .A3(new_n725_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n730_), .A2(new_n731_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n488_), .B1(new_n772_), .B2(KEYINPUT113), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n747_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n768_), .B1(new_n775_), .B2(new_n751_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n752_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n548_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(KEYINPUT57), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n607_), .B1(new_n779_), .B2(new_n762_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT118), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(new_n607_), .C1(new_n779_), .C2(new_n762_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n717_), .A3(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n765_), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n767_), .A2(new_n428_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G113gat), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n429_), .A2(G113gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n766_), .B2(new_n789_), .ZN(G1340gat));
  NAND3_X1  g589(.A1(new_n767_), .A2(new_n502_), .A3(new_n786_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G120gat), .ZN(new_n792_));
  INV_X1    g591(.A(G120gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n639_), .B2(KEYINPUT60), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(KEYINPUT60), .B2(new_n793_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n766_), .B2(new_n795_), .ZN(G1341gat));
  INV_X1    g595(.A(new_n766_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G127gat), .B1(new_n797_), .B2(new_n539_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n767_), .A2(new_n786_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n538_), .A2(G127gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT119), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n798_), .B1(new_n799_), .B2(new_n801_), .ZN(G1342gat));
  XNOR2_X1  g601(.A(KEYINPUT121), .B(G134gat), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n602_), .A2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT122), .ZN(new_n805_));
  INV_X1    g604(.A(G134gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n766_), .B2(new_n547_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT120), .B(new_n806_), .C1(new_n766_), .C2(new_n547_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n799_), .A2(new_n805_), .B1(new_n809_), .B2(new_n810_), .ZN(G1343gat));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n778_), .B2(KEYINPUT57), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n757_), .A2(new_n761_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n753_), .A2(KEYINPUT116), .A3(new_n754_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n538_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n716_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n375_), .A2(new_n404_), .A3(new_n543_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n818_), .A2(new_n619_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n428_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n502_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g623(.A1(new_n820_), .A2(new_n539_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT61), .B(G155gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1346gat));
  INV_X1    g626(.A(G162gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n820_), .A2(new_n828_), .A3(new_n548_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n820_), .A2(new_n602_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1347gat));
  INV_X1    g630(.A(KEYINPUT22), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n618_), .A2(new_n289_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n586_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n784_), .A2(new_n832_), .A3(new_n428_), .A4(new_n834_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n835_), .A2(KEYINPUT62), .A3(new_n211_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n784_), .A2(new_n834_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n429_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n211_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(KEYINPUT62), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n836_), .B1(new_n840_), .B2(new_n841_), .ZN(G1348gat));
  INV_X1    g641(.A(new_n837_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G176gat), .B1(new_n843_), .B2(new_n502_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n833_), .A2(new_n639_), .A3(new_n212_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT123), .B1(new_n764_), .B2(new_n376_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n818_), .A2(new_n847_), .A3(new_n375_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT124), .B(new_n845_), .C1(new_n846_), .C2(new_n848_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n844_), .B1(new_n851_), .B2(new_n852_), .ZN(G1349gat));
  NOR3_X1   g652(.A1(new_n837_), .A2(new_n316_), .A3(new_n817_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n833_), .A2(new_n607_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n847_), .B1(new_n818_), .B2(new_n375_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n756_), .A2(new_n762_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n538_), .B1(new_n857_), .B2(new_n815_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT123), .B(new_n376_), .C1(new_n858_), .C2(new_n716_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n855_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G183gat), .B1(new_n860_), .B2(KEYINPUT125), .ZN(new_n861_));
  INV_X1    g660(.A(new_n855_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n854_), .B1(new_n861_), .B2(new_n865_), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n837_), .B2(new_n524_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n548_), .A2(new_n317_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n837_), .B2(new_n868_), .ZN(G1351gat));
  NAND3_X1  g668(.A1(new_n375_), .A2(new_n404_), .A3(new_n288_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT126), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n870_), .A2(KEYINPUT126), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n619_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n818_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n428_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n502_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n877_), .B(new_n878_), .Z(G1353gat));
  NAND2_X1  g678(.A1(new_n874_), .A2(new_n538_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n880_), .B2(new_n881_), .ZN(G1354gat));
  INV_X1    g683(.A(G218gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n874_), .A2(new_n885_), .A3(new_n548_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n818_), .A2(new_n524_), .A3(new_n873_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1355gat));
endmodule


