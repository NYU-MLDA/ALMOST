//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_,
    new_n995_;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203_));
  INV_X1    g002(.A(G29gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G36gat), .ZN(new_n205_));
  INV_X1    g004(.A(G36gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G29gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(G29gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(G36gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT72), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217_));
  INV_X1    g016(.A(G1gat), .ZN(new_n218_));
  INV_X1    g017(.A(G8gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G1gat), .B(G8gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n216_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n223_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n216_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n225_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n215_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n213_), .A3(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n226_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  OAI22_X1  g033(.A1(new_n224_), .A2(new_n225_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n202_), .B1(new_n237_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n240_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n235_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n202_), .A3(new_n241_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G85gat), .B(G92gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT6), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(G99gat), .A3(G106gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  AOI211_X1 g058(.A(KEYINPUT8), .B(new_n250_), .C1(new_n254_), .C2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT8), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT7), .ZN(new_n262_));
  INV_X1    g061(.A(G99gat), .ZN(new_n263_));
  INV_X1    g062(.A(G106gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n257_), .B1(G99gat), .B2(G106gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n255_), .A2(KEYINPUT6), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n251_), .B(new_n265_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n250_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n261_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n264_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT64), .ZN(new_n274_));
  AND2_X1   g073(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n264_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT9), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n281_), .A2(G85gat), .A3(G92gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G85gat), .A2(G92gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n281_), .A2(KEYINPUT65), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n281_), .A2(KEYINPUT65), .ZN(new_n286_));
  OAI22_X1  g085(.A1(new_n282_), .A2(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n288_));
  INV_X1    g087(.A(G85gat), .ZN(new_n289_));
  INV_X1    g088(.A(G92gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT9), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n283_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n292_), .A3(new_n259_), .ZN(new_n293_));
  OAI22_X1  g092(.A1(new_n260_), .A2(new_n270_), .B1(new_n280_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT66), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n274_), .A2(new_n279_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n288_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n283_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n297_), .A2(new_n298_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n299_), .A3(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n300_), .B(new_n301_), .C1(new_n270_), .C2(new_n260_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G57gat), .B(G64gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n305_));
  XOR2_X1   g104(.A(G71gat), .B(G78gat), .Z(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT12), .B1(new_n303_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n310_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n295_), .A2(new_n312_), .A3(new_n302_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n294_), .A2(KEYINPUT12), .A3(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G230gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n311_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n302_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n268_), .A2(new_n269_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT8), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n268_), .A2(new_n261_), .A3(new_n269_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n301_), .B1(new_n323_), .B2(new_n300_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n310_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n303_), .A2(KEYINPUT68), .A3(new_n310_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n313_), .A2(KEYINPUT67), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n295_), .A2(new_n330_), .A3(new_n312_), .A4(new_n302_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .A4(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n318_), .B1(new_n317_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G120gat), .B(G148gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT5), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G176gat), .B(G204gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT70), .B1(new_n333_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n333_), .B2(KEYINPUT69), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n329_), .A2(new_n331_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT68), .B1(new_n303_), .B2(new_n310_), .ZN(new_n342_));
  AOI211_X1 g141(.A(new_n326_), .B(new_n312_), .C1(new_n295_), .C2(new_n302_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n316_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n318_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n339_), .B1(new_n340_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT13), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n346_), .B1(new_n345_), .B2(new_n318_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n332_), .A2(new_n317_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n318_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(KEYINPUT69), .A3(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n350_), .A2(KEYINPUT70), .A3(new_n353_), .A4(new_n337_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n348_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n349_), .B1(new_n348_), .B2(new_n354_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n249_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(new_n352_), .A3(new_n338_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n351_), .A2(new_n352_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n338_), .B1(new_n361_), .B2(new_n346_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n362_), .B2(new_n353_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n354_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT13), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n348_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT71), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n248_), .B1(new_n357_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G113gat), .B(G120gat), .Z(new_n374_));
  NOR2_X1   g173(.A1(new_n374_), .A2(KEYINPUT83), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n375_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(KEYINPUT83), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n377_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT94), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT2), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n395_));
  NOR3_X1   g194(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n394_), .B(new_n395_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(KEYINPUT3), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n390_), .B(new_n391_), .C1(new_n398_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n392_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(new_n399_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n388_), .A2(new_n389_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n391_), .B(KEYINPUT1), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n385_), .A2(new_n386_), .A3(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n406_), .A2(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n401_), .A2(KEYINPUT3), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n396_), .A2(new_n397_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n391_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n406_), .A2(new_n415_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n411_), .A2(new_n405_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n379_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n382_), .A2(new_n383_), .A3(new_n381_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT94), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n410_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n376_), .B(KEYINPUT83), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(new_n381_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n427_), .B2(new_n409_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n426_), .ZN(new_n430_));
  AND4_X1   g229(.A1(new_n423_), .A2(new_n429_), .A3(new_n430_), .A4(new_n409_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n422_), .B(KEYINPUT4), .C1(new_n428_), .C2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n409_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT95), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n432_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n422_), .B(new_n435_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n373_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n386_), .B1(new_n385_), .B2(new_n409_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n417_), .A2(new_n420_), .A3(KEYINPUT94), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n429_), .A2(new_n430_), .A3(new_n409_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT93), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n427_), .A2(new_n423_), .A3(new_n409_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n444_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n437_), .B1(new_n448_), .B2(KEYINPUT4), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(new_n373_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT101), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n372_), .B1(new_n448_), .B2(new_n435_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT101), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n439_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n441_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT103), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G78gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G228gat), .A2(G233gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(G197gat), .B(G204gat), .Z(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT21), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G197gat), .B(G204gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT21), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G211gat), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n466_), .A2(G218gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT89), .B1(new_n466_), .B2(G218gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n461_), .B(KEYINPUT21), .C1(new_n467_), .C2(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(KEYINPUT90), .A3(new_n471_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n459_), .A2(new_n460_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT29), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n472_), .ZN(new_n479_));
  OAI211_X1 g278(.A(G228gat), .B(G233gat), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n458_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n476_), .A2(new_n480_), .A3(new_n458_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(G106gat), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n483_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n264_), .B1(new_n485_), .B2(new_n481_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT91), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n484_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n417_), .A2(new_n477_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT28), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G22gat), .B(G50gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n489_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(KEYINPUT91), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n474_), .A2(new_n475_), .ZN(new_n500_));
  INV_X1    g299(.A(G169gat), .ZN(new_n501_));
  INV_X1    g300(.A(G176gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(KEYINPUT81), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(KEYINPUT81), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G183gat), .A2(G190gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT23), .ZN(new_n509_));
  NOR3_X1   g308(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT26), .B(G190gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT80), .B(G183gat), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT25), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n514_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n508_), .B(KEYINPUT23), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(G190gat), .B2(new_n515_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n501_), .B2(KEYINPUT22), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G169gat), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n502_), .B(new_n523_), .C1(new_n524_), .C2(new_n522_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n521_), .B(new_n525_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n500_), .A2(new_n519_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n528_));
  INV_X1    g327(.A(new_n509_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(new_n505_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT25), .B(G183gat), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n510_), .B1(new_n513_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n509_), .B1(G183gat), .B2(G190gat), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n503_), .B1(new_n524_), .B2(new_n502_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n530_), .A2(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n528_), .B1(new_n536_), .B2(new_n472_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n527_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G226gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT19), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G8gat), .B(G36gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G64gat), .B(G92gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n526_), .B1(new_n512_), .B2(new_n518_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n540_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n528_), .B1(new_n535_), .B2(new_n479_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n541_), .A2(new_n546_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n546_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n551_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n549_), .B1(new_n527_), .B2(new_n537_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT27), .B1(new_n552_), .B2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n552_), .A2(KEYINPUT27), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n548_), .A2(new_n550_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n540_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n540_), .B2(new_n538_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n553_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n557_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G71gat), .B(G99gat), .ZN(new_n564_));
  INV_X1    g363(.A(G43gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n547_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(G15gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT30), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n567_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(KEYINPUT85), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n427_), .B(KEYINPUT31), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(KEYINPUT85), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n457_), .A2(new_n499_), .A3(new_n563_), .A4(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n441_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n454_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n453_), .B1(new_n452_), .B2(new_n439_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n541_), .A2(new_n551_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n546_), .A2(KEYINPUT32), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT100), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n554_), .A2(new_n555_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n584_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n586_), .A2(new_n589_), .B1(new_n561_), .B2(new_n585_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n582_), .A2(new_n590_), .A3(KEYINPUT102), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT102), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n561_), .A2(new_n585_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n583_), .A2(KEYINPUT100), .A3(new_n585_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n588_), .B1(new_n587_), .B2(new_n584_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n455_), .B2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n434_), .A2(new_n435_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n432_), .A2(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT99), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(KEYINPUT99), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n373_), .B1(new_n448_), .B2(new_n436_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n552_), .A2(new_n556_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n449_), .A2(new_n450_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n605_), .B2(KEYINPUT33), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n452_), .A2(new_n439_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT98), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n611_));
  AOI211_X1 g410(.A(new_n611_), .B(new_n608_), .C1(new_n452_), .C2(new_n439_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n603_), .B(new_n606_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n591_), .A2(new_n597_), .A3(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n496_), .A2(new_n498_), .A3(new_n563_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n614_), .A2(new_n499_), .B1(new_n457_), .B2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n578_), .B1(new_n616_), .B2(new_n577_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n368_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT76), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n231_), .A2(new_n233_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT34), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI22_X1  g423(.A1(new_n620_), .A2(new_n294_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n295_), .A2(new_n302_), .A3(new_n216_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(KEYINPUT74), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n624_), .A2(new_n621_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n625_), .B(new_n626_), .C1(KEYINPUT74), .C2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT36), .Z(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(KEYINPUT36), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n630_), .A2(new_n632_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n619_), .B1(new_n641_), .B2(KEYINPUT37), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT75), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  INV_X1    g444(.A(new_n637_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT75), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n644_), .A2(new_n645_), .A3(new_n640_), .A4(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n633_), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n651_), .A2(new_n639_), .B1(new_n647_), .B2(KEYINPUT75), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n652_), .A2(new_n619_), .A3(new_n645_), .A4(new_n644_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(G127gat), .B(G155gat), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT16), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G183gat), .B(G211gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(G231gat), .A2(G233gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n223_), .B(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n310_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n226_), .A2(new_n659_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n223_), .B1(G231gat), .B2(G233gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n312_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n658_), .B1(new_n665_), .B2(KEYINPUT17), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n658_), .A2(KEYINPUT17), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n665_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(KEYINPUT77), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(KEYINPUT77), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n654_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n618_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT104), .ZN(new_n676_));
  INV_X1    g475(.A(new_n457_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n618_), .A2(new_n678_), .A3(new_n674_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n676_), .A2(new_n218_), .A3(new_n677_), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT38), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n652_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n644_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n617_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n673_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n368_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G1gat), .B1(new_n689_), .B2(new_n457_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n680_), .A2(new_n681_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n690_), .A3(new_n691_), .ZN(G1324gat));
  NOR2_X1   g491(.A1(new_n563_), .A2(G8gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n676_), .A2(new_n679_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n676_), .A2(KEYINPUT105), .A3(new_n679_), .A4(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G8gat), .B1(new_n689_), .B2(new_n563_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT39), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n700_), .A3(KEYINPUT40), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1325gat));
  INV_X1    g504(.A(new_n577_), .ZN(new_n706_));
  OR3_X1    g505(.A1(new_n675_), .A2(G15gat), .A3(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n689_), .A2(new_n706_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT41), .B1(new_n708_), .B2(G15gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT106), .B(new_n707_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1326gat));
  OAI21_X1  g514(.A(G22gat), .B1(new_n689_), .B2(new_n499_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT42), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n499_), .A2(G22gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT107), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n675_), .B2(new_n719_), .ZN(G1327gat));
  AND2_X1   g519(.A1(new_n368_), .A2(new_n673_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n617_), .A2(new_n722_), .A3(new_n654_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n617_), .B2(new_n654_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT44), .B(new_n721_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n727_), .A2(G29gat), .A3(new_n677_), .A4(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n686_), .A2(new_n688_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n618_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n204_), .B1(new_n731_), .B2(new_n457_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n729_), .A2(new_n732_), .ZN(G1328gat));
  NOR2_X1   g532(.A1(new_n563_), .A2(G36gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n618_), .A2(new_n730_), .A3(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n736_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n618_), .A2(new_n730_), .A3(new_n738_), .A4(new_n734_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n563_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n727_), .A2(new_n741_), .A3(new_n728_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n742_), .B2(G36gat), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n745_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n743_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1329gat));
  NAND4_X1  g549(.A1(new_n727_), .A2(G43gat), .A3(new_n577_), .A4(new_n728_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n565_), .B1(new_n731_), .B2(new_n706_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(G1330gat));
  INV_X1    g554(.A(new_n499_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n727_), .A2(G50gat), .A3(new_n756_), .A4(new_n728_), .ZN(new_n757_));
  INV_X1    g556(.A(G50gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n731_), .B2(new_n499_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1331gat));
  NAND2_X1  g559(.A1(new_n357_), .A2(new_n367_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n762_), .A2(new_n248_), .A3(new_n617_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n674_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n677_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n687_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n247_), .A2(new_n673_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n769_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n768_), .A2(new_n457_), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n766_), .B2(new_n771_), .ZN(G1332gat));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n773_), .A3(new_n741_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n768_), .A2(new_n563_), .A3(new_n770_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(G64gat), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n776_), .A2(KEYINPUT48), .A3(new_n773_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n774_), .B1(new_n778_), .B2(new_n779_), .ZN(G1333gat));
  INV_X1    g579(.A(G71gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n765_), .A2(new_n781_), .A3(new_n577_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n768_), .A2(new_n706_), .A3(new_n770_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(G71gat), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n784_), .A2(KEYINPUT49), .A3(new_n781_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n756_), .A2(new_n458_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT113), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n765_), .A2(new_n790_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n768_), .A2(new_n499_), .A3(new_n770_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(G78gat), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G78gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n795_), .B2(new_n796_), .ZN(G1335gat));
  NAND2_X1  g596(.A1(new_n763_), .A2(new_n730_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n289_), .B1(new_n798_), .B2(new_n457_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT114), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n357_), .A2(new_n367_), .A3(new_n673_), .A4(new_n248_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n617_), .A2(new_n654_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT43), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n617_), .A2(new_n722_), .A3(new_n654_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n806_), .A2(new_n289_), .A3(new_n457_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n800_), .A2(new_n807_), .ZN(G1336gat));
  OAI21_X1  g607(.A(G92gat), .B1(new_n806_), .B2(new_n563_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n798_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n290_), .A3(new_n741_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1337gat));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n277_), .A3(new_n577_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n805_), .A2(new_n577_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n814_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT115), .B1(new_n814_), .B2(G99gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n813_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT51), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n813_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1338gat));
  NOR2_X1   g620(.A1(new_n499_), .A2(G106gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n810_), .A2(KEYINPUT116), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824_));
  INV_X1    g623(.A(new_n822_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n798_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n805_), .A2(KEYINPUT117), .A3(new_n756_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n801_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n756_), .B(new_n829_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n828_), .A2(new_n832_), .A3(KEYINPUT52), .A4(G106gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n827_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n830_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n264_), .B1(new_n835_), .B2(KEYINPUT117), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(new_n836_), .B2(new_n832_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT53), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n828_), .A2(G106gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n832_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n833_), .A4(new_n827_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n838_), .A2(new_n844_), .ZN(G1339gat));
  AND3_X1   g644(.A1(new_n650_), .A2(new_n653_), .A3(new_n769_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT118), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n846_), .A2(new_n365_), .A3(new_n366_), .A4(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(KEYINPUT54), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n847_), .A2(KEYINPUT118), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n225_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n227_), .A2(new_n855_), .ZN(new_n856_));
  OAI221_X1 g655(.A(new_n244_), .B1(new_n856_), .B2(new_n234_), .C1(new_n224_), .C2(new_n855_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n245_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n348_), .A2(new_n354_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n348_), .A2(KEYINPUT119), .A3(new_n354_), .A4(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n247_), .A2(new_n358_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n311_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n315_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n317_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n318_), .B1(new_n868_), .B2(KEYINPUT55), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n867_), .A2(new_n870_), .A3(new_n317_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n337_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT56), .B(new_n337_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n864_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n863_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(KEYINPUT57), .A3(new_n686_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n876_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n685_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n358_), .A2(new_n858_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n884_), .A2(KEYINPUT58), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n654_), .B1(new_n884_), .B2(KEYINPUT58), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n879_), .A2(new_n882_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n854_), .B1(new_n888_), .B2(new_n673_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n577_), .A2(new_n499_), .A3(new_n563_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n457_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(G113gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n247_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n885_), .A2(new_n886_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n685_), .B1(new_n863_), .B2(new_n877_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(KEYINPUT57), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n688_), .B1(new_n900_), .B2(new_n882_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT59), .B(new_n891_), .C1(new_n901_), .C2(new_n854_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n248_), .B1(new_n897_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n895_), .B1(new_n903_), .B2(new_n894_), .ZN(G1340gat));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905_));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n897_), .A2(new_n902_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n762_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n893_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n761_), .B2(KEYINPUT60), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(KEYINPUT60), .B2(new_n906_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n905_), .B1(new_n908_), .B2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n761_), .B1(new_n897_), .B2(new_n902_), .ZN(new_n914_));
  OAI221_X1 g713(.A(KEYINPUT121), .B1(new_n909_), .B2(new_n911_), .C1(new_n914_), .C2(new_n906_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1341gat));
  INV_X1    g715(.A(G127gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n893_), .A2(new_n917_), .A3(new_n688_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n673_), .B1(new_n897_), .B2(new_n902_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n917_), .ZN(G1342gat));
  INV_X1    g719(.A(G134gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n893_), .A2(new_n921_), .A3(new_n685_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n654_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n897_), .B2(new_n902_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n924_), .B2(new_n921_), .ZN(G1343gat));
  NOR2_X1   g724(.A1(new_n889_), .A2(new_n577_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n677_), .A3(new_n615_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n248_), .ZN(new_n928_));
  INV_X1    g727(.A(G141gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1344gat));
  NOR2_X1   g729(.A1(new_n927_), .A2(new_n761_), .ZN(new_n931_));
  INV_X1    g730(.A(G148gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1345gat));
  NOR2_X1   g732(.A1(new_n927_), .A2(new_n673_), .ZN(new_n934_));
  XOR2_X1   g733(.A(KEYINPUT61), .B(G155gat), .Z(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1346gat));
  OAI21_X1  g735(.A(G162gat), .B1(new_n927_), .B2(new_n923_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n686_), .A2(G162gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n927_), .B2(new_n938_), .ZN(G1347gat));
  NAND2_X1  g738(.A1(new_n888_), .A2(new_n673_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n854_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n457_), .A2(new_n741_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n943_), .A2(new_n756_), .A3(new_n706_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n942_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(KEYINPUT124), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n942_), .A2(new_n944_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n946_), .A2(new_n949_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n247_), .A2(new_n524_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n247_), .B(new_n944_), .C1(new_n901_), .C2(new_n854_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n942_), .A2(KEYINPUT122), .A3(new_n247_), .A4(new_n944_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n958_));
  OAI21_X1  g757(.A(G169gat), .B1(new_n958_), .B2(KEYINPUT123), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  AOI22_X1  g759(.A1(new_n957_), .A2(new_n960_), .B1(KEYINPUT123), .B2(new_n958_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n958_), .A2(KEYINPUT123), .ZN(new_n962_));
  AOI211_X1 g761(.A(new_n962_), .B(new_n959_), .C1(new_n955_), .C2(new_n956_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n952_), .B1(new_n961_), .B2(new_n963_), .ZN(G1348gat));
  NAND3_X1  g763(.A1(new_n950_), .A2(new_n502_), .A3(new_n762_), .ZN(new_n965_));
  OAI21_X1  g764(.A(G176gat), .B1(new_n947_), .B2(new_n761_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1349gat));
  AOI21_X1  g766(.A(new_n515_), .B1(new_n945_), .B2(new_n688_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n673_), .A2(new_n531_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n950_), .B2(new_n969_), .ZN(G1350gat));
  NOR2_X1   g769(.A1(new_n686_), .A2(new_n514_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n950_), .A2(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(G190gat), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n923_), .B1(new_n946_), .B2(new_n949_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n972_), .B1(new_n973_), .B2(new_n974_), .ZN(G1351gat));
  NOR2_X1   g774(.A1(new_n943_), .A2(new_n499_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n942_), .A2(new_n706_), .A3(new_n976_), .ZN(new_n977_));
  INV_X1    g776(.A(new_n977_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(new_n247_), .ZN(new_n979_));
  XNOR2_X1  g778(.A(new_n979_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g779(.A1(new_n978_), .A2(new_n762_), .ZN(new_n981_));
  AND2_X1   g780(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n982_));
  NOR2_X1   g781(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n981_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n984_), .B1(new_n981_), .B2(new_n982_), .ZN(G1353gat));
  OAI22_X1  g784(.A1(new_n977_), .A2(new_n673_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987_));
  XNOR2_X1  g786(.A(KEYINPUT63), .B(G211gat), .ZN(new_n988_));
  NAND4_X1  g787(.A1(new_n926_), .A2(new_n688_), .A3(new_n976_), .A4(new_n988_), .ZN(new_n989_));
  AND3_X1   g788(.A1(new_n986_), .A2(new_n987_), .A3(new_n989_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n987_), .B1(new_n986_), .B2(new_n989_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(new_n990_), .A2(new_n991_), .ZN(G1354gat));
  XOR2_X1   g791(.A(KEYINPUT127), .B(G218gat), .Z(new_n993_));
  NOR3_X1   g792(.A1(new_n977_), .A2(new_n923_), .A3(new_n993_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n978_), .A2(new_n685_), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n994_), .B1(new_n995_), .B2(new_n993_), .ZN(G1355gat));
endmodule


