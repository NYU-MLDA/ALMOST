//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  OAI211_X1 g000(.A(G85gat), .B(G92gat), .C1(KEYINPUT65), .C2(KEYINPUT9), .ZN(new_n202_));
  OAI211_X1 g001(.A(KEYINPUT65), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT10), .B(G99gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G106gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n204_), .A2(new_n207_), .A3(new_n212_), .ZN(new_n213_));
  OR3_X1    g012(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT66), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n212_), .A2(new_n214_), .A3(new_n216_), .A4(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G85gat), .B(G92gat), .Z(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT8), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n223_), .A3(new_n220_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n213_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G29gat), .B(G36gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(KEYINPUT73), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(KEYINPUT73), .ZN(new_n228_));
  XOR2_X1   g027(.A(G43gat), .B(G50gat), .Z(new_n229_));
  OR3_X1    g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n229_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n225_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n225_), .A2(KEYINPUT75), .A3(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G232gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT34), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT35), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT74), .B(KEYINPUT15), .Z(new_n241_));
  NAND3_X1  g040(.A1(new_n230_), .A2(new_n231_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n241_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n213_), .A2(KEYINPUT69), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n222_), .A2(new_n224_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n204_), .A2(new_n207_), .A3(new_n212_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n240_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n237_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n239_), .A2(KEYINPUT35), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n237_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT76), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G190gat), .B(G218gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G134gat), .B(G162gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT36), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n256_), .A2(KEYINPUT76), .A3(new_n257_), .A4(new_n262_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n261_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT36), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n271_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G64gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G57gat), .ZN(new_n281_));
  INV_X1    g080(.A(G57gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G64gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n283_), .A3(KEYINPUT11), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT68), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT11), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n282_), .A2(G64gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n280_), .A2(G57gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(G71gat), .A2(G78gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G71gat), .A2(G78gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n290_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT11), .B1(new_n281_), .B2(new_n283_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G71gat), .B(G78gat), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n299_), .A2(KEYINPUT67), .A3(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n289_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT67), .B1(new_n299_), .B2(new_n300_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n297_), .B(new_n290_), .C1(new_n286_), .C2(KEYINPUT11), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n303_), .A2(new_n285_), .A3(new_n288_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n251_), .A2(KEYINPUT12), .A3(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n219_), .A2(new_n223_), .A3(new_n220_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n223_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n248_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(new_n306_), .ZN(new_n311_));
  AND2_X1   g110(.A1(G230gat), .A2(G233gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n306_), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n314_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  AOI211_X1 g117(.A(KEYINPUT71), .B(new_n316_), .C1(new_n310_), .C2(new_n306_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n307_), .B(new_n313_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n247_), .A2(new_n248_), .B1(new_n305_), .B2(new_n302_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n311_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G120gat), .B(G148gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT5), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G176gat), .B(G204gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n323_), .B(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G231gat), .A2(G233gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n306_), .B(new_n335_), .Z(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT78), .B(G15gat), .ZN(new_n337_));
  INV_X1    g136(.A(G22gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G1gat), .ZN(new_n340_));
  INV_X1    g139(.A(G8gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT14), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G8gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT79), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n344_), .B(KEYINPUT79), .Z(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n342_), .A3(new_n339_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n336_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G155gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G183gat), .B(G211gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT17), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(KEYINPUT17), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n350_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT81), .B1(new_n350_), .B2(new_n356_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(new_n358_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n279_), .A2(new_n334_), .A3(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT87), .B(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT31), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT88), .ZN(new_n368_));
  INV_X1    g167(.A(G15gat), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n370_), .A2(new_n371_), .A3(G227gat), .A4(G233gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(KEYINPUT84), .A2(KEYINPUT26), .ZN(new_n377_));
  NAND2_X1  g176(.A1(KEYINPUT84), .A2(KEYINPUT26), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(G190gat), .A3(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT25), .B(G183gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT83), .B(G190gat), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n379_), .B(new_n380_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G183gat), .A3(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT23), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n386_), .B2(KEYINPUT23), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n395_), .B2(KEYINPUT24), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n383_), .A2(new_n390_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n386_), .A2(KEYINPUT23), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n385_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n382_), .B2(G183gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT86), .ZN(new_n401_));
  INV_X1    g200(.A(G169gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT22), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G176gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT22), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(KEYINPUT86), .A3(G169gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n400_), .A2(new_n392_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n397_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT30), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n376_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n409_), .B(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n375_), .A3(new_n374_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G127gat), .B(G134gat), .Z(new_n415_));
  XOR2_X1   g214(.A(G113gat), .B(G120gat), .Z(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n411_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n366_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n411_), .A2(new_n414_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n417_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n365_), .A3(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n431_));
  INV_X1    g230(.A(G141gat), .ZN(new_n432_));
  INV_X1    g231(.A(G148gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n432_), .A2(new_n433_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n430_), .B(new_n434_), .C1(new_n435_), .C2(KEYINPUT2), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT90), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n439_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n429_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G141gat), .B(G148gat), .Z(new_n443_));
  NAND3_X1  g242(.A1(new_n428_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G155gat), .A3(G162gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n446_), .A3(new_n427_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT89), .B1(new_n428_), .B2(KEYINPUT1), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n443_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n442_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n442_), .A2(KEYINPUT91), .A3(new_n449_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n417_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n417_), .A2(new_n450_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G225gat), .A2(G233gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT101), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n454_), .A2(KEYINPUT4), .A3(new_n455_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT102), .B(KEYINPUT4), .Z(new_n466_));
  NAND4_X1  g265(.A1(new_n452_), .A2(new_n453_), .A3(new_n417_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n457_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n459_), .B(new_n464_), .C1(new_n465_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n454_), .A2(new_n455_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n457_), .B(new_n467_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n464_), .B1(new_n473_), .B2(new_n459_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n426_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G226gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT19), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G211gat), .B(G218gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G197gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G204gat), .ZN(new_n484_));
  INV_X1    g283(.A(G204gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G197gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n487_), .A3(KEYINPUT95), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT95), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n486_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(new_n481_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n480_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n484_), .A2(new_n486_), .A3(KEYINPUT92), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT21), .B1(new_n484_), .B2(KEYINPUT92), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT21), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n485_), .A2(G197gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n484_), .A2(new_n486_), .A3(KEYINPUT92), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(KEYINPUT93), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n492_), .A2(new_n503_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n487_), .A2(new_n479_), .A3(new_n497_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT20), .B1(new_n507_), .B2(new_n409_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n492_), .B2(new_n503_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(G183gat), .A2(G190gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n390_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT22), .B(G169gat), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n393_), .B1(new_n513_), .B2(new_n404_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G190gat), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n395_), .A2(new_n515_), .B1(new_n380_), .B2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n518_));
  AOI22_X1  g317(.A1(new_n518_), .A2(new_n394_), .B1(new_n385_), .B2(new_n398_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n512_), .A2(new_n514_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n509_), .A2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n478_), .B1(new_n508_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT100), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n504_), .A2(new_n520_), .A3(new_n506_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n478_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n397_), .A2(new_n408_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT20), .B1(new_n509_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n523_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT20), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n507_), .B2(new_n409_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n478_), .B1(new_n509_), .B2(new_n520_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT100), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G8gat), .B(G36gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT18), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G64gat), .B(G92gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n522_), .A2(new_n529_), .A3(new_n533_), .A4(new_n538_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT27), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n541_), .A2(KEYINPUT27), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT97), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n507_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n509_), .A2(KEYINPUT97), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n520_), .A2(KEYINPUT104), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n520_), .A2(KEYINPUT104), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n525_), .B1(new_n551_), .B2(new_n531_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n508_), .A2(new_n478_), .A3(new_n521_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n539_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n545_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n544_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n452_), .A2(KEYINPUT29), .A3(new_n453_), .ZN(new_n558_));
  INV_X1    g357(.A(G228gat), .ZN(new_n559_));
  INV_X1    g358(.A(G233gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n558_), .A2(new_n507_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n450_), .B2(KEYINPUT29), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n566_));
  AOI211_X1 g365(.A(KEYINPUT96), .B(new_n566_), .C1(new_n442_), .C2(new_n449_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n509_), .A2(KEYINPUT97), .ZN(new_n569_));
  AOI211_X1 g368(.A(new_n546_), .B(new_n505_), .C1(new_n492_), .C2(new_n503_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n563_), .B1(new_n571_), .B2(new_n561_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G78gat), .B(G106gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n557_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n452_), .A2(new_n453_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n566_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G22gat), .B(G50gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT28), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n577_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n561_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n563_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n582_), .A2(new_n574_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n574_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n585_));
  OAI22_X1  g384(.A1(new_n575_), .A2(new_n581_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n573_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n572_), .A2(new_n574_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n557_), .A3(new_n589_), .A4(new_n580_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n476_), .A2(new_n556_), .A3(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n586_), .A2(new_n590_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n464_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n467_), .A2(new_n458_), .ZN(new_n595_));
  OAI221_X1 g394(.A(new_n594_), .B1(new_n471_), .B2(new_n458_), .C1(new_n465_), .C2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n540_), .A2(new_n541_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n469_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n538_), .A2(KEYINPUT32), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n522_), .A2(new_n529_), .A3(new_n533_), .A4(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n551_), .A2(new_n531_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n553_), .B1(new_n602_), .B2(new_n478_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n601_), .B1(new_n603_), .B2(new_n600_), .ZN(new_n604_));
  OAI22_X1  g403(.A1(new_n597_), .A2(new_n599_), .B1(new_n604_), .B2(new_n475_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n593_), .A2(new_n605_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n543_), .A2(new_n542_), .B1(new_n545_), .B2(new_n554_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n591_), .A3(new_n475_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n426_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n592_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  OR2_X1    g413(.A1(new_n349_), .A2(new_n232_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n349_), .A2(new_n232_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n244_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n621_), .A2(new_n348_), .A3(new_n346_), .A4(new_n242_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n349_), .B2(new_n232_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT82), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n614_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n617_), .A2(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n614_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n628_), .A2(KEYINPUT82), .A3(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n363_), .A2(new_n611_), .A3(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n475_), .B(KEYINPUT105), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n340_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n273_), .B(KEYINPUT106), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n611_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n334_), .A2(new_n631_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n362_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n475_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n635_), .A2(new_n636_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n637_), .A2(new_n645_), .A3(new_n646_), .ZN(G1324gat));
  OAI21_X1  g446(.A(G8gat), .B1(new_n644_), .B2(new_n607_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT39), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n633_), .A2(new_n341_), .A3(new_n556_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n644_), .B2(new_n610_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT41), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n633_), .A2(new_n369_), .A3(new_n426_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n644_), .B2(new_n593_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n633_), .A2(new_n338_), .A3(new_n591_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n274_), .B1(new_n266_), .B2(new_n272_), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n271_), .B(new_n275_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n426_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n664_), .B(new_n667_), .C1(new_n668_), .C2(new_n592_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT109), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n556_), .A2(new_n591_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n475_), .A3(new_n426_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n475_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n674_));
  AOI22_X1  g473(.A1(new_n605_), .A2(new_n593_), .B1(new_n674_), .B2(new_n607_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n675_), .B2(new_n426_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n664_), .A4(new_n667_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n611_), .B2(new_n279_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n670_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n641_), .A2(new_n362_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n634_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G29gat), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n362_), .A2(new_n277_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n676_), .A2(new_n631_), .A3(new_n334_), .A4(new_n689_), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n690_), .A2(G29gat), .A3(new_n475_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1328gat));
  NOR3_X1   g491(.A1(new_n690_), .A2(G36gat), .A3(new_n607_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT45), .Z(new_n694_));
  AND3_X1   g493(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n681_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT44), .B1(new_n680_), .B2(new_n681_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT110), .B1(new_n697_), .B2(new_n556_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n684_), .A2(KEYINPUT110), .A3(new_n556_), .A4(new_n685_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n694_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT46), .B(new_n694_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n697_), .A2(new_n706_), .A3(G43gat), .A4(new_n426_), .ZN(new_n707_));
  INV_X1    g506(.A(G43gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n686_), .A2(new_n708_), .A3(new_n610_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n690_), .A2(new_n610_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT111), .B1(new_n710_), .B2(new_n708_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT47), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n707_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1330gat));
  OAI21_X1  g515(.A(G50gat), .B1(new_n686_), .B2(new_n593_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n593_), .A2(G50gat), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT112), .Z(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n690_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(new_n334_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n640_), .A2(new_n632_), .A3(new_n721_), .A4(new_n362_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(new_n282_), .A3(new_n475_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n611_), .A2(new_n631_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n667_), .A2(new_n642_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n721_), .A3(new_n725_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT113), .Z(new_n727_));
  AOI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n634_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n728_), .A2(KEYINPUT114), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(KEYINPUT114), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n723_), .B1(new_n729_), .B2(new_n730_), .ZN(G1332gat));
  OAI21_X1  g530(.A(G64gat), .B1(new_n722_), .B2(new_n607_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT48), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n280_), .A3(new_n556_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n722_), .B2(new_n610_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n738_), .A3(new_n426_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n722_), .B2(new_n593_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n593_), .A2(G78gat), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT115), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n727_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1335gat));
  INV_X1    g545(.A(G85gat), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n334_), .A2(new_n362_), .A3(new_n631_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n680_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n749_), .B2(new_n673_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n724_), .A2(new_n721_), .A3(new_n689_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n751_), .A2(G85gat), .A3(new_n687_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1336gat));
  INV_X1    g552(.A(G92gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n749_), .B2(new_n556_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n751_), .A2(G92gat), .A3(new_n607_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1337gat));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n751_), .A2(new_n610_), .A3(new_n205_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n749_), .A2(new_n426_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G99gat), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762_));
  AND4_X1   g561(.A1(new_n758_), .A2(new_n761_), .A3(new_n762_), .A4(KEYINPUT51), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n762_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT51), .B1(new_n761_), .B2(new_n758_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1338gat));
  OR3_X1    g565(.A1(new_n751_), .A2(new_n593_), .A3(new_n206_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n749_), .A2(new_n591_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n767_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  NAND3_X1  g575(.A1(new_n320_), .A2(new_n322_), .A3(new_n328_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n631_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n311_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n307_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n312_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n320_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT71), .B1(new_n321_), .B2(new_n316_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n315_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n307_), .A4(new_n313_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n781_), .A2(new_n783_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n327_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n327_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n778_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n622_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n619_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n629_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n622_), .A2(new_n623_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n618_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n614_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n329_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n277_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT57), .B(new_n277_), .C1(new_n793_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n796_), .A2(new_n799_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n777_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(new_n777_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n792_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n791_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n789_), .A2(new_n810_), .A3(new_n790_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n667_), .B1(new_n814_), .B2(KEYINPUT58), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n807_), .A2(new_n808_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n327_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n810_), .B2(new_n792_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n813_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n803_), .B(new_n804_), .C1(new_n815_), .C2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n642_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT54), .B1(new_n363_), .B2(new_n631_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n725_), .A2(new_n826_), .A3(new_n632_), .A4(new_n334_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n824_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n671_), .A2(new_n426_), .A3(new_n634_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n823_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n820_), .A2(new_n821_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n814_), .A2(KEYINPUT58), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n667_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(KEYINPUT120), .A3(new_n803_), .A4(new_n804_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n835_), .A2(new_n642_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n828_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n831_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n833_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n632_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n847_), .A3(new_n631_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n845_), .B2(new_n334_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n334_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n843_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(G1341gat));
  NAND2_X1  g653(.A1(new_n362_), .A2(G127gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT122), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n833_), .B(new_n856_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G127gat), .B1(new_n843_), .B2(new_n362_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1342gat));
  OAI21_X1  g659(.A(G134gat), .B1(new_n845_), .B2(new_n279_), .ZN(new_n861_));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n843_), .A2(new_n862_), .A3(new_n639_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n426_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n687_), .A2(new_n593_), .A3(new_n556_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n362_), .B1(new_n823_), .B2(new_n834_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n828_), .B1(new_n869_), .B2(new_n839_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n867_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n870_), .A2(KEYINPUT123), .A3(new_n426_), .A4(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n631_), .B1(new_n868_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G141gat), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n432_), .B(new_n631_), .C1(new_n868_), .C2(new_n872_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1344gat));
  OAI21_X1  g675(.A(new_n721_), .B1(new_n868_), .B2(new_n872_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G148gat), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n433_), .B(new_n721_), .C1(new_n868_), .C2(new_n872_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1345gat));
  OAI21_X1  g679(.A(new_n362_), .B1(new_n868_), .B2(new_n872_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n882_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n362_), .B(new_n884_), .C1(new_n868_), .C2(new_n872_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1346gat));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n887_), .B(new_n639_), .C1(new_n868_), .C2(new_n872_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n866_), .A2(new_n867_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT123), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n866_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n279_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n888_), .B1(new_n892_), .B2(new_n887_), .ZN(G1347gat));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n607_), .A2(new_n610_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n687_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n591_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n632_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n824_), .B2(new_n828_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n402_), .B1(new_n900_), .B2(KEYINPUT124), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(new_n899_), .C1(new_n824_), .C2(new_n828_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n894_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  INV_X1    g704(.A(new_n900_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n905_), .B1(new_n513_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(G169gat), .A3(new_n903_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT125), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n901_), .A2(new_n894_), .A3(new_n903_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(KEYINPUT62), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n912_), .ZN(G1348gat));
  NAND2_X1  g712(.A1(new_n830_), .A2(new_n897_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n404_), .B1(new_n914_), .B2(new_n334_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n842_), .A2(new_n593_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n896_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(new_n721_), .A3(G176gat), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n915_), .B(new_n916_), .C1(new_n917_), .C2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n829_), .A2(new_n898_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G176gat), .B1(new_n921_), .B2(new_n721_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n917_), .A2(new_n919_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT126), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n924_), .ZN(G1349gat));
  NOR3_X1   g724(.A1(new_n914_), .A2(new_n380_), .A3(new_n642_), .ZN(new_n926_));
  INV_X1    g725(.A(G183gat), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n842_), .A2(new_n593_), .A3(new_n362_), .A4(new_n918_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n914_), .B2(new_n279_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n921_), .A2(new_n516_), .A3(new_n639_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1351gat));
  NAND2_X1  g731(.A1(new_n674_), .A2(new_n556_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n866_), .A2(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n632_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(new_n483_), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n334_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n485_), .ZN(G1353gat));
  AOI21_X1  g738(.A(new_n642_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n866_), .A2(new_n934_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT127), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n941_), .B(new_n943_), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n935_), .B2(new_n279_), .ZN(new_n945_));
  OR2_X1    g744(.A1(new_n638_), .A2(G218gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n935_), .B2(new_n946_), .ZN(G1355gat));
endmodule


