//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(KEYINPUT78), .A2(G1gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT78), .A2(G1gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(G8gat), .A3(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(KEYINPUT79), .A3(KEYINPUT14), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT79), .B1(new_n208_), .B2(KEYINPUT14), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n205_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(G1gat), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(KEYINPUT14), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n209_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n218_), .B2(new_n205_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n204_), .B1(new_n213_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT73), .B(G29gat), .ZN(new_n221_));
  INV_X1    g020(.A(G36gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G43gat), .B(G50gat), .Z(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n221_), .B(G36gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(new_n224_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n212_), .A2(G1gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n218_), .A2(new_n214_), .A3(new_n205_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(G8gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n220_), .A2(new_n230_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n230_), .B1(new_n220_), .B2(new_n233_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n203_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n220_), .A2(new_n233_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n229_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT15), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n227_), .A2(new_n224_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n223_), .A2(new_n225_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT15), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n220_), .A2(new_n245_), .A3(new_n233_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n246_), .A3(new_n202_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n237_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249_));
  INV_X1    g048(.A(G169gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G197gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n248_), .A2(KEYINPUT80), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n248_), .B2(KEYINPUT80), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT19), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT90), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT21), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT88), .B(G197gat), .ZN(new_n263_));
  INV_X1    g062(.A(G204gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n252_), .B2(new_n264_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n252_), .A2(G204gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n263_), .B2(G204gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n268_), .A2(new_n269_), .B1(new_n262_), .B2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G211gat), .B(G218gat), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n271_), .A2(new_n274_), .A3(new_n262_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT23), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(G183gat), .B2(G190gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT22), .B(G169gat), .ZN(new_n284_));
  INV_X1    g083(.A(G176gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G190gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n289_));
  AND2_X1   g088(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n250_), .A2(new_n285_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT24), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT24), .A3(new_n282_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n291_), .A2(new_n280_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n287_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n278_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n276_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT91), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n281_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n281_), .A2(new_n299_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n286_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(new_n295_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n298_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n261_), .B1(new_n297_), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT18), .B(G64gat), .ZN(new_n306_));
  INV_X1    g105(.A(G92gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n278_), .A2(new_n296_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n259_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n298_), .A2(new_n303_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n311_), .A2(KEYINPUT20), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n305_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n310_), .B1(new_n305_), .B2(new_n314_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318_));
  INV_X1    g117(.A(G141gat), .ZN(new_n319_));
  INV_X1    g118(.A(G148gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n321_), .A2(new_n323_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(G141gat), .B2(G148gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT85), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n327_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n332_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341_));
  INV_X1    g140(.A(G113gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G120gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(G120gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n343_), .B(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n339_), .A3(new_n332_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(KEYINPUT4), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n350_), .A3(new_n344_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n345_), .A2(new_n352_), .A3(new_n348_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT0), .B(G57gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G85gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(G1gat), .B(G29gat), .Z(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT92), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  OR3_X1    g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n349_), .A2(new_n352_), .A3(new_n351_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n345_), .A2(new_n348_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT93), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n359_), .B(new_n367_), .C1(new_n369_), .C2(new_n352_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n363_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n317_), .A2(new_n366_), .A3(new_n370_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n354_), .A2(new_n355_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n359_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n361_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n310_), .A2(KEYINPUT32), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n305_), .A2(new_n314_), .A3(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n297_), .A2(new_n304_), .A3(new_n261_), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n381_));
  NAND3_X1  g180(.A1(new_n311_), .A2(new_n313_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n259_), .B2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n377_), .B(new_n379_), .C1(new_n383_), .C2(new_n378_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n371_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n315_), .A2(new_n316_), .A3(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n386_), .A2(KEYINPUT94), .A3(new_n370_), .A4(new_n366_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n374_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G227gat), .A2(G233gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(KEYINPUT30), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n296_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G15gat), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT83), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G71gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G99gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n396_), .A2(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n389_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT84), .A3(new_n399_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n347_), .B(KEYINPUT31), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n389_), .B(new_n405_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT87), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n278_), .A2(new_n410_), .B1(G228gat), .B2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT28), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n278_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n415_), .A2(KEYINPUT28), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(KEYINPUT28), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(new_n278_), .A3(new_n421_), .A4(new_n417_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n419_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n414_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n427_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n413_), .A3(new_n425_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n388_), .A2(new_n409_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n310_), .B(KEYINPUT96), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n383_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n315_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n317_), .A2(KEYINPUT27), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n377_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n409_), .A2(new_n430_), .A3(new_n428_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n409_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n438_), .B(new_n439_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n432_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT74), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT7), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT7), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT67), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  AOI211_X1 g249(.A(G99gat), .B(G106gat), .C1(new_n446_), .C2(KEYINPUT7), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT68), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n447_), .A2(new_n445_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n457_), .B(new_n458_), .C1(new_n459_), .C2(new_n445_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n452_), .A2(new_n456_), .A3(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT8), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n458_), .B1(new_n459_), .B2(new_n445_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(new_n455_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n464_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n463_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT9), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT9), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n463_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n462_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT65), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G99gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT10), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT10), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G99gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(G106gat), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n455_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n475_), .A2(KEYINPUT65), .A3(new_n462_), .A4(new_n477_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n480_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT66), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n480_), .A2(new_n490_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n467_), .A2(new_n472_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT15), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT15), .B1(new_n242_), .B2(new_n243_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n444_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n489_), .A2(new_n491_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n468_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n471_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n245_), .B(KEYINPUT74), .C1(new_n497_), .C2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n497_), .A2(new_n499_), .A3(new_n230_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G232gat), .A2(G233gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT71), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n502_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n505_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n508_), .A2(new_n505_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G190gat), .B(G218gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G134gat), .ZN(new_n515_));
  INV_X1    g314(.A(G162gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT76), .Z(new_n520_));
  AND3_X1   g319(.A1(new_n509_), .A2(new_n513_), .A3(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n517_), .B(KEYINPUT36), .Z(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n521_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT77), .ZN(new_n526_));
  AND4_X1   g325(.A1(new_n511_), .A2(new_n501_), .A3(new_n512_), .A4(new_n503_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n511_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n509_), .A2(KEYINPUT77), .A3(new_n513_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n522_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n521_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n525_), .B1(new_n534_), .B2(new_n524_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n238_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(KEYINPUT11), .ZN(new_n538_));
  INV_X1    g337(.A(G57gat), .ZN(new_n539_));
  INV_X1    g338(.A(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G57gat), .A2(G64gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n538_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546_));
  INV_X1    g345(.A(G71gat), .ZN(new_n547_));
  INV_X1    g346(.A(G78gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT69), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(KEYINPUT69), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n544_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(new_n543_), .A3(new_n551_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n537_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT16), .B(G183gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G211gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT17), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n537_), .A2(new_n557_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n558_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n558_), .A2(new_n564_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n557_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n554_), .A2(new_n556_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n489_), .A2(new_n491_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n571_), .B(new_n572_), .C1(new_n498_), .C2(new_n471_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(KEYINPUT12), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n575_), .B(new_n557_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n264_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(G176gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n578_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n589_), .B2(new_n580_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n587_), .A2(KEYINPUT70), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT70), .B1(new_n587_), .B2(new_n590_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT13), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT70), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n586_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n589_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n587_), .A2(KEYINPUT70), .A3(new_n590_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n569_), .A2(new_n593_), .A3(new_n600_), .ZN(new_n601_));
  AND4_X1   g400(.A1(new_n257_), .A2(new_n443_), .A3(new_n535_), .A4(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n206_), .A2(new_n207_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n377_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT38), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT13), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n598_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n256_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT97), .ZN(new_n611_));
  INV_X1    g410(.A(new_n569_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n432_), .B2(new_n442_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n534_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT98), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n439_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n605_), .B1(new_n619_), .B2(new_n214_), .ZN(G1324gat));
  INV_X1    g419(.A(new_n438_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n602_), .A2(new_n204_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n621_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(G8gat), .ZN(new_n625_));
  AOI211_X1 g424(.A(KEYINPUT39), .B(new_n204_), .C1(new_n615_), .C2(new_n621_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g427(.A(new_n409_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n629_));
  INV_X1    g428(.A(G15gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT99), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n409_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n618_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n611_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(G15gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n631_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n602_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n631_), .A2(new_n637_), .A3(KEYINPUT41), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(G1326gat));
  AOI21_X1  g442(.A(new_n431_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n644_));
  INV_X1    g443(.A(G22gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT100), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n431_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(G22gat), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n602_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n650_), .A3(KEYINPUT42), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(G1327gat));
  AOI21_X1  g455(.A(new_n535_), .B1(new_n432_), .B2(new_n442_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n610_), .B(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n659_), .A2(KEYINPUT44), .A3(new_n661_), .A4(new_n612_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n534_), .A2(new_n524_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n525_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n658_), .B1(new_n443_), .B2(new_n665_), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT43), .B(new_n535_), .C1(new_n432_), .C2(new_n442_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n661_), .B(new_n612_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n662_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n377_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(KEYINPUT101), .A3(new_n377_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(G29gat), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n534_), .B1(new_n432_), .B2(new_n442_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n679_), .A2(G29gat), .A3(new_n439_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n682_), .A2(KEYINPUT102), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n662_), .A2(new_n670_), .A3(new_n621_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(KEYINPUT102), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n677_), .A2(new_n222_), .A3(new_n610_), .A4(new_n612_), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n687_), .A2(KEYINPUT45), .A3(new_n438_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT45), .B1(new_n687_), .B2(new_n438_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AND4_X1   g489(.A1(new_n683_), .A2(new_n685_), .A3(new_n686_), .A4(new_n690_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n684_), .A2(G36gat), .B1(new_n689_), .B2(new_n688_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n683_), .B1(new_n692_), .B2(new_n686_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1329gat));
  NAND3_X1  g493(.A1(new_n671_), .A2(G43gat), .A3(new_n632_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G43gat), .B1(new_n678_), .B2(new_n632_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT103), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT47), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n700_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1330gat));
  NAND2_X1  g501(.A1(new_n671_), .A2(new_n647_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G50gat), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n431_), .A2(G50gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n679_), .B2(new_n705_), .ZN(G1331gat));
  NAND4_X1  g505(.A1(new_n613_), .A2(new_n609_), .A3(new_n256_), .A4(new_n535_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT104), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n377_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n614_), .A2(new_n608_), .A3(new_n257_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(new_n377_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(G57gat), .B2(new_n711_), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n540_), .B1(new_n710_), .B2(new_n621_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT48), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n621_), .A2(new_n540_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT105), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n708_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1333gat));
  AOI21_X1  g517(.A(new_n547_), .B1(new_n710_), .B2(new_n632_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT49), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n708_), .A2(new_n547_), .A3(new_n632_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1334gat));
  AOI21_X1  g521(.A(new_n548_), .B1(new_n710_), .B2(new_n647_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT50), .Z(new_n724_));
  NAND2_X1  g523(.A1(new_n647_), .A2(new_n548_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT106), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n708_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(G1335gat));
  NOR3_X1   g527(.A1(new_n608_), .A2(new_n257_), .A3(new_n569_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n677_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT107), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n377_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n659_), .A2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n377_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n732_), .B1(new_n735_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g535(.A(G92gat), .B1(new_n731_), .B2(new_n621_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n438_), .A2(new_n307_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n733_), .B2(new_n738_), .ZN(G1337gat));
  NAND2_X1  g538(.A1(new_n482_), .A2(new_n484_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n731_), .A2(new_n740_), .A3(new_n632_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n659_), .A2(new_n632_), .A3(new_n729_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G99gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT108), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(new_n743_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(KEYINPUT51), .A3(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1338gat));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n659_), .A2(new_n753_), .A3(new_n647_), .A4(new_n729_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n647_), .B(new_n729_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT110), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(new_n756_), .A3(G106gat), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(G106gat), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n730_), .A2(KEYINPUT107), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n730_), .A2(KEYINPUT107), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n761_), .B(new_n647_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT109), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n731_), .A2(new_n766_), .A3(new_n761_), .A4(new_n647_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n754_), .A2(new_n756_), .A3(G106gat), .A4(new_n758_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n760_), .A2(new_n768_), .A3(new_n771_), .A4(new_n769_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1339gat));
  OAI21_X1  g574(.A(new_n587_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n574_), .A2(new_n588_), .A3(new_n576_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n579_), .A2(KEYINPUT55), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n589_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n779_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n777_), .B1(new_n783_), .B2(new_n586_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n781_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT55), .B(new_n588_), .C1(new_n574_), .C2(new_n576_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n778_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n776_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n253_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n202_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n239_), .A2(new_n246_), .A3(new_n203_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n253_), .B1(new_n237_), .B2(new_n247_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT113), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n246_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n796_), .A2(new_n236_), .A3(new_n202_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n203_), .B1(new_n239_), .B2(new_n234_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n253_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n796_), .A2(new_n236_), .A3(new_n203_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n202_), .B1(new_n239_), .B2(new_n234_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n790_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AND4_X1   g603(.A1(new_n599_), .A2(new_n597_), .A3(new_n795_), .A4(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n534_), .B1(new_n789_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI221_X1 g607(.A(new_n534_), .B1(KEYINPUT114), .B2(KEYINPUT57), .C1(new_n789_), .C2(new_n805_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n795_), .A2(new_n804_), .A3(new_n587_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n585_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n810_), .B(KEYINPUT58), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n665_), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n809_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n612_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n608_), .A2(new_n535_), .A3(new_n256_), .A4(new_n569_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n601_), .A2(KEYINPUT54), .A3(new_n256_), .A4(new_n535_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(new_n377_), .A3(new_n438_), .A4(new_n441_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n257_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n621_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT115), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n831_), .A2(new_n377_), .A3(new_n441_), .A4(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n256_), .B1(new_n830_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n828_), .B1(new_n835_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g635(.A(new_n830_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n834_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n609_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT116), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n841_), .B(new_n609_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(G120gat), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n346_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n827_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n346_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n827_), .A2(new_n847_), .A3(new_n569_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n612_), .B1(new_n830_), .B2(new_n834_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT117), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n852_), .B(new_n848_), .C1(new_n849_), .C2(new_n847_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1342gat));
  INV_X1    g653(.A(new_n534_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G134gat), .B1(new_n827_), .B2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT118), .B(G134gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n830_), .B2(new_n834_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n858_), .B2(new_n665_), .ZN(G1343gat));
  AND3_X1   g658(.A1(new_n831_), .A2(new_n377_), .A3(new_n440_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n257_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT119), .B(G141gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n609_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n569_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  AOI21_X1  g667(.A(G162gat), .B1(new_n860_), .B2(new_n855_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n535_), .A2(new_n516_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n860_), .B2(new_n870_), .ZN(G1347gat));
  AOI211_X1 g670(.A(new_n377_), .B(new_n438_), .C1(new_n819_), .C2(new_n824_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n872_), .A2(new_n441_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n257_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n441_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT120), .B1(new_n876_), .B2(new_n256_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(G169gat), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n873_), .A2(new_n257_), .A3(new_n284_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n875_), .A2(KEYINPUT62), .A3(new_n877_), .A4(G169gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n876_), .A2(new_n608_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n285_), .ZN(G1349gat));
  AOI21_X1  g684(.A(new_n290_), .B1(KEYINPUT121), .B2(new_n289_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n873_), .A2(new_n569_), .A3(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(G183gat), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT121), .B(new_n888_), .C1(new_n876_), .C2(new_n612_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1350gat));
  NAND3_X1  g691(.A1(new_n873_), .A2(new_n288_), .A3(new_n855_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G190gat), .B1(new_n876_), .B2(new_n535_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  AND2_X1   g694(.A1(new_n872_), .A2(new_n440_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G197gat), .B1(new_n896_), .B2(new_n257_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n872_), .A2(new_n440_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n900_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n901_), .A2(KEYINPUT123), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(KEYINPUT123), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n898_), .A2(new_n899_), .B1(new_n902_), .B2(new_n903_), .ZN(G1352gat));
  NOR2_X1   g703(.A1(new_n900_), .A2(new_n608_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT125), .B(G204gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1353gat));
  NOR2_X1   g706(.A1(new_n900_), .A2(new_n612_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT63), .B(G211gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n908_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT126), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n910_), .B(new_n914_), .C1(new_n908_), .C2(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1354gat));
  AOI21_X1  g715(.A(G218gat), .B1(new_n896_), .B2(new_n855_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n665_), .A2(G218gat), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT127), .Z(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n896_), .B2(new_n919_), .ZN(G1355gat));
endmodule


