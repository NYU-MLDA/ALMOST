//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT87), .Z(new_n208_));
  OR2_X1    g007(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n210_));
  INV_X1    g009(.A(G155gat), .ZN(new_n211_));
  INV_X1    g010(.A(G162gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n209_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n205_), .B1(new_n208_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n206_), .A3(new_n214_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT89), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT90), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n202_), .A2(KEYINPUT88), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT3), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT3), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n204_), .B(KEYINPUT2), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n220_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n220_), .B1(new_n219_), .B2(new_n225_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n217_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT28), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n219_), .A2(new_n225_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT90), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n216_), .B1(new_n232_), .B2(new_n226_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G22gat), .B(G50gat), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n230_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n230_), .B2(new_n236_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G78gat), .B(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT96), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n245_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n229_), .A2(KEYINPUT96), .A3(KEYINPUT29), .ZN(new_n247_));
  XOR2_X1   g046(.A(G211gat), .B(G218gat), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT94), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT94), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n249_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n253_), .B(KEYINPUT94), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n250_), .B(new_n251_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n246_), .A2(new_n247_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT93), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(G228gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(G228gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(KEYINPUT95), .ZN(new_n268_));
  INV_X1    g067(.A(new_n252_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n250_), .A2(new_n251_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n255_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n253_), .A2(new_n254_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n269_), .B(new_n270_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT95), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n256_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n268_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(new_n266_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT92), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n233_), .A2(new_n278_), .A3(new_n235_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT92), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n277_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n244_), .B1(new_n267_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT97), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n267_), .A2(new_n244_), .A3(new_n281_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AOI211_X1 g084(.A(KEYINPUT97), .B(new_n244_), .C1(new_n267_), .C2(new_n281_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n242_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n282_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n284_), .A3(new_n240_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT23), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT81), .B(G190gat), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n291_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G169gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(KEYINPUT26), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n305_));
  OR3_X1    g104(.A1(new_n305_), .A2(new_n292_), .A3(KEYINPUT26), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n292_), .B2(KEYINPUT26), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n303_), .A2(new_n304_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(G183gat), .B2(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT84), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n295_), .A2(KEYINPUT84), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n294_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(G176gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT83), .ZN(new_n321_));
  OR3_X1    g120(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT83), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n317_), .B(new_n323_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n302_), .B1(new_n315_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G71gat), .B(G99gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G43gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n326_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n330_), .B(G15gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT30), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT31), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n329_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G127gat), .B(G134gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n336_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT0), .B(G57gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n229_), .A2(new_n341_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n233_), .A2(new_n342_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT4), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n229_), .A2(new_n356_), .A3(new_n341_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n353_), .A2(KEYINPUT99), .A3(new_n355_), .A4(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n355_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT99), .B1(new_n362_), .B2(new_n353_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n350_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT99), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT4), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(new_n361_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n367_), .A2(new_n349_), .A3(new_n359_), .A4(new_n358_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n345_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n273_), .A2(new_n274_), .A3(new_n256_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n274_), .B1(new_n273_), .B2(new_n256_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n376_), .B2(new_n326_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n304_), .A2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n296_), .A2(new_n322_), .A3(new_n320_), .A4(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n301_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n314_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT98), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n310_), .A2(new_n311_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n295_), .A2(KEYINPUT84), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n293_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n301_), .B1(new_n389_), .B2(new_n383_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT98), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n381_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n259_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n373_), .B1(new_n377_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n373_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT20), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n376_), .B2(new_n326_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n394_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT18), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n396_), .A2(new_n406_), .A3(new_n401_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT27), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT102), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n396_), .A2(new_n401_), .A3(KEYINPUT102), .A4(new_n406_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n326_), .A2(new_n268_), .A3(new_n275_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n394_), .A2(new_n390_), .A3(new_n380_), .ZN(new_n419_));
  XOR2_X1   g218(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n373_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT101), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n382_), .B1(new_n298_), .B2(new_n296_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n308_), .A2(new_n314_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n325_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n424_), .B1(new_n276_), .B2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n429_), .B(new_n397_), .C1(new_n394_), .C2(new_n393_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT101), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n431_), .B(new_n373_), .C1(new_n418_), .C2(new_n421_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n423_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n416_), .B1(new_n433_), .B2(new_n407_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT103), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n415_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n415_), .B2(new_n434_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n411_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n290_), .A2(new_n371_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n289_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n284_), .A2(new_n283_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n288_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n286_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n440_), .B1(new_n444_), .B2(new_n242_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n368_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n368_), .A2(new_n446_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n353_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n351_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n350_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n408_), .B(new_n409_), .C1(new_n449_), .C2(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n447_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n402_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n454_), .B2(new_n433_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n369_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n445_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n415_), .A2(new_n434_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT103), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n415_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n410_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(new_n290_), .A3(new_n370_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n345_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n439_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G113gat), .B(G141gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT80), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G169gat), .B(G197gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n473_));
  INV_X1    g272(.A(G8gat), .ZN(new_n474_));
  INV_X1    g273(.A(G1gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT72), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT72), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(G1gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n473_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT72), .B(G1gat), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n482_), .C2(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G15gat), .B(G22gat), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT74), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT74), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n489_), .A3(new_n486_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n489_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n494_));
  AOI211_X1 g293(.A(KEYINPUT74), .B(new_n485_), .C1(new_n481_), .C2(new_n483_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497_));
  XOR2_X1   g296(.A(G29gat), .B(G36gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT68), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G29gat), .B(G36gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n503_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n497_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(KEYINPUT15), .A3(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n492_), .A2(new_n496_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n492_), .A2(new_n496_), .A3(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT79), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n505_), .A2(new_n506_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n472_), .B(new_n512_), .C1(new_n514_), .C2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n491_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n494_), .A2(new_n495_), .A3(new_n493_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n515_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n492_), .A2(new_n496_), .A3(new_n516_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n492_), .A2(new_n496_), .A3(KEYINPUT78), .A4(new_n516_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n472_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n471_), .B1(new_n519_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n472_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n492_), .A2(new_n496_), .A3(new_n516_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n530_), .A2(new_n517_), .A3(KEYINPUT78), .ZN(new_n531_));
  INV_X1    g330(.A(new_n526_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n518_), .A3(new_n470_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n466_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G127gat), .B(G155gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G183gat), .B(G211gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT75), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n492_), .A2(new_n496_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n547_));
  INV_X1    g346(.A(G64gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G57gat), .ZN(new_n549_));
  INV_X1    g348(.A(G57gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(G64gat), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n549_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT11), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n551_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT66), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT11), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(KEYINPUT11), .B(new_n561_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n546_), .A2(new_n547_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n565_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT17), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n543_), .B1(new_n568_), .B2(new_n541_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT77), .B1(new_n566_), .B2(new_n567_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n576_));
  INV_X1    g375(.A(G99gat), .ZN(new_n577_));
  INV_X1    g376(.A(G106gat), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT6), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT6), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(G99gat), .A3(G106gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G85gat), .ZN(new_n583_));
  INV_X1    g382(.A(G92gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT9), .A3(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n578_), .A3(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n586_), .A2(KEYINPUT9), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n582_), .A2(new_n587_), .A3(new_n590_), .A4(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n586_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT64), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n594_), .B(new_n595_), .C1(G99gat), .C2(G106gat), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n577_), .B(new_n578_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n593_), .B1(new_n598_), .B2(new_n582_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n592_), .B1(new_n599_), .B2(KEYINPUT8), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n593_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(KEYINPUT65), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT65), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n596_), .A2(new_n597_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n582_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT8), .B(new_n602_), .C1(new_n604_), .C2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n601_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n510_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT35), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n614_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n515_), .A2(new_n601_), .A3(new_n608_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n610_), .A2(new_n616_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n617_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n507_), .A2(new_n509_), .B1(new_n601_), .B2(new_n608_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n615_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n576_), .B1(new_n623_), .B2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n619_), .A2(new_n622_), .A3(KEYINPUT69), .A4(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n626_), .B(KEYINPUT36), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n623_), .A2(new_n632_), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT70), .B(new_n575_), .C1(new_n631_), .C2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT70), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(new_n633_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n636_), .B2(KEYINPUT37), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT71), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n623_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n619_), .A2(new_n622_), .A3(KEYINPUT71), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n640_), .A3(new_n632_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n631_), .A2(new_n575_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n634_), .B1(new_n637_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT67), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT5), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n565_), .A2(new_n601_), .A3(new_n608_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n602_), .A2(KEYINPUT8), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n606_), .A2(new_n582_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n603_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n564_), .B(new_n563_), .C1(new_n655_), .C2(new_n600_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n656_), .A3(KEYINPUT12), .ZN(new_n657_));
  INV_X1    g456(.A(new_n565_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT12), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n609_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n651_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n650_), .B1(new_n652_), .B2(new_n656_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n649_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n649_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n645_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(KEYINPUT67), .A3(new_n663_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT13), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n574_), .A2(new_n644_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n536_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(new_n482_), .A3(new_n369_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(KEYINPUT38), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT104), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n631_), .A2(new_n641_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n466_), .A2(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n574_), .A2(new_n535_), .A3(new_n671_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n475_), .B1(new_n683_), .B2(new_n369_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n675_), .B2(KEYINPUT38), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n677_), .A2(new_n685_), .ZN(G1324gat));
  NAND3_X1  g485(.A1(new_n674_), .A2(new_n474_), .A3(new_n438_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n474_), .B1(new_n683_), .B2(new_n438_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT39), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n688_), .A2(new_n689_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1325gat));
  OAI21_X1  g494(.A(G15gat), .B1(new_n682_), .B2(new_n465_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT41), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n673_), .A2(G15gat), .A3(new_n465_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n682_), .B2(new_n445_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n445_), .A2(G22gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n673_), .B2(new_n702_), .ZN(G1327gat));
  NOR3_X1   g502(.A1(new_n671_), .A2(new_n573_), .A3(new_n678_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n536_), .A2(new_n704_), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n705_), .A2(G29gat), .A3(new_n370_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n671_), .A2(new_n535_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n574_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n445_), .A2(new_n438_), .A3(new_n369_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n452_), .B1(new_n446_), .B2(new_n368_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n448_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n712_), .A2(new_n713_), .B1(new_n369_), .B2(new_n456_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n290_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n465_), .B1(new_n711_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n439_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n710_), .B1(new_n718_), .B2(new_n644_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n345_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n710_), .B(new_n644_), .C1(new_n720_), .C2(new_n439_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n709_), .C1(new_n719_), .C2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n466_), .B2(new_n643_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n708_), .B1(new_n724_), .B2(new_n721_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n723_), .B(new_n369_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n727_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT106), .B1(new_n727_), .B2(G29gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n706_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT107), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(new_n706_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1328gat));
  NOR3_X1   g533(.A1(new_n705_), .A2(G36gat), .A3(new_n462_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT45), .Z(new_n736_));
  INV_X1    g535(.A(G36gat), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n725_), .A2(new_n726_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n739_), .B(new_n708_), .C1(new_n724_), .C2(new_n721_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n738_), .A2(new_n740_), .A3(new_n462_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n736_), .B(KEYINPUT46), .C1(new_n737_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1329gat));
  NOR2_X1   g545(.A1(new_n738_), .A2(new_n740_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(G43gat), .A3(new_n345_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n705_), .A2(new_n465_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(G43gat), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g550(.A1(new_n705_), .A2(G50gat), .A3(new_n445_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n723_), .B(new_n290_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G50gat), .B1(new_n753_), .B2(new_n754_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT109), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n752_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1331gat));
  INV_X1    g560(.A(new_n535_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n466_), .A2(new_n762_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n574_), .A2(new_n644_), .A3(new_n670_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n550_), .B1(new_n765_), .B2(new_n370_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n670_), .A2(new_n762_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n574_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n680_), .A2(new_n769_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n770_), .A2(new_n550_), .A3(new_n370_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n766_), .B1(new_n771_), .B2(KEYINPUT110), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(KEYINPUT110), .B2(new_n771_), .ZN(G1332gat));
  INV_X1    g572(.A(new_n770_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n548_), .B1(new_n774_), .B2(new_n438_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT48), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n775_), .A2(new_n776_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n438_), .A2(new_n548_), .ZN(new_n780_));
  OAI22_X1  g579(.A1(new_n778_), .A2(new_n779_), .B1(new_n765_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(G1333gat));
  OAI21_X1  g582(.A(G71gat), .B1(new_n770_), .B2(new_n465_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT49), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n465_), .A2(G71gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n765_), .B2(new_n786_), .ZN(G1334gat));
  OAI21_X1  g586(.A(G78gat), .B1(new_n770_), .B2(new_n445_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT50), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n445_), .A2(G78gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n765_), .B2(new_n790_), .ZN(G1335gat));
  NOR3_X1   g590(.A1(new_n573_), .A2(new_n678_), .A3(new_n670_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n763_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n583_), .A3(new_n369_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n724_), .A2(new_n721_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n768_), .A2(new_n573_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(new_n369_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n799_), .B2(new_n583_), .ZN(G1336gat));
  NOR3_X1   g599(.A1(new_n793_), .A2(G92gat), .A3(new_n462_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n438_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(G92gat), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT112), .Z(G1337gat));
  AOI21_X1  g603(.A(new_n577_), .B1(new_n798_), .B2(new_n345_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n345_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n794_), .B2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n796_), .A2(new_n290_), .A3(new_n797_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(G106gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT114), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(new_n813_), .A3(G106gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(KEYINPUT52), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n794_), .A2(new_n578_), .A3(new_n290_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n812_), .B2(KEYINPUT52), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT53), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n812_), .A2(KEYINPUT52), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n815_), .A4(new_n817_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(G1339gat));
  NAND2_X1  g622(.A1(new_n657_), .A2(new_n660_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n650_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n661_), .A2(KEYINPUT55), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n657_), .A2(new_n651_), .A3(new_n660_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT115), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n657_), .A2(new_n831_), .A3(new_n651_), .A4(new_n660_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n827_), .A2(new_n828_), .A3(new_n830_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n649_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT56), .ZN(new_n835_));
  INV_X1    g634(.A(new_n649_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n830_), .A2(new_n832_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT55), .B1(new_n824_), .B2(new_n650_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n826_), .B(new_n651_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n836_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n835_), .A2(new_n843_), .A3(new_n667_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n512_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n472_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n847_), .B2(new_n846_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n531_), .A2(new_n532_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n471_), .B1(new_n850_), .B2(new_n472_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n533_), .A2(new_n518_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n849_), .A2(new_n851_), .B1(new_n852_), .B2(new_n471_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n844_), .A2(new_n845_), .A3(KEYINPUT58), .A4(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n665_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n853_), .A2(new_n855_), .A3(KEYINPUT58), .A4(new_n835_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT119), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n853_), .A2(new_n855_), .A3(new_n835_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n643_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n665_), .B1(new_n528_), .B2(new_n534_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n842_), .B1(new_n841_), .B2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n834_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n867_), .A2(KEYINPUT117), .B1(new_n669_), .B2(new_n853_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n863_), .A2(new_n865_), .A3(new_n869_), .A4(new_n866_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n679_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n862_), .B1(new_n871_), .B2(KEYINPUT57), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n867_), .A2(KEYINPUT117), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n853_), .A2(new_n669_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n870_), .A3(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT57), .A3(new_n678_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n574_), .B1(new_n872_), .B2(new_n877_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n573_), .A2(new_n643_), .A3(new_n535_), .A4(new_n670_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n290_), .A2(new_n438_), .A3(new_n465_), .A4(new_n370_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G113gat), .B1(new_n885_), .B2(new_n762_), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(KEYINPUT120), .Z(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n884_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT59), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n762_), .A2(G113gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n887_), .B1(new_n890_), .B2(new_n891_), .ZN(G1340gat));
  INV_X1    g691(.A(G120gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n670_), .B2(KEYINPUT60), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n885_), .B(new_n894_), .C1(KEYINPUT60), .C2(new_n893_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT121), .Z(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT122), .B1(new_n889_), .B2(new_n670_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G120gat), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n889_), .A2(KEYINPUT122), .A3(new_n670_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1341gat));
  OAI21_X1  g699(.A(G127gat), .B1(new_n889_), .B2(new_n574_), .ZN(new_n901_));
  OR3_X1    g700(.A1(new_n888_), .A2(G127gat), .A3(new_n574_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1342gat));
  AOI21_X1  g702(.A(G134gat), .B1(new_n885_), .B2(new_n679_), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT123), .Z(new_n905_));
  AND2_X1   g704(.A1(new_n644_), .A2(G134gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n890_), .B2(new_n906_), .ZN(G1343gat));
  NAND2_X1  g706(.A1(new_n875_), .A2(new_n678_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n910_), .A2(new_n876_), .A3(new_n862_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n881_), .B1(new_n911_), .B2(new_n574_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n345_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n445_), .A2(new_n438_), .A3(new_n370_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n762_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n671_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g719(.A1(new_n915_), .A2(new_n574_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT61), .B(G155gat), .Z(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n915_), .B2(new_n643_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n679_), .A2(new_n212_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n915_), .B2(new_n925_), .ZN(G1347gat));
  NOR3_X1   g725(.A1(new_n462_), .A2(new_n371_), .A3(new_n290_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n912_), .A2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n318_), .B1(new_n929_), .B2(new_n762_), .ZN(new_n930_));
  XOR2_X1   g729(.A(new_n930_), .B(KEYINPUT62), .Z(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT124), .B1(new_n912_), .B2(new_n928_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933_));
  AOI22_X1  g732(.A1(new_n908_), .A2(new_n909_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n573_), .B1(new_n934_), .B2(new_n876_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n933_), .B(new_n927_), .C1(new_n935_), .C2(new_n881_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n938_));
  AND2_X1   g737(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n937_), .B(new_n762_), .C1(new_n938_), .C2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n931_), .A2(new_n940_), .ZN(G1348gat));
  NAND3_X1  g740(.A1(new_n937_), .A2(new_n319_), .A3(new_n671_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n912_), .A2(new_n670_), .A3(new_n928_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n319_), .B2(new_n943_), .ZN(G1349gat));
  AOI21_X1  g743(.A(G183gat), .B1(new_n929_), .B2(new_n573_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n574_), .A2(new_n304_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n937_), .B2(new_n946_), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n937_), .A2(new_n378_), .A3(new_n679_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n933_), .B1(new_n883_), .B2(new_n927_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n912_), .A2(KEYINPUT124), .A3(new_n928_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n644_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n949_), .B1(new_n952_), .B2(G190gat), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n643_), .B1(new_n932_), .B2(new_n936_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n954_), .A2(KEYINPUT125), .A3(new_n292_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n948_), .B1(new_n953_), .B2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  OAI211_X1 g757(.A(KEYINPUT126), .B(new_n948_), .C1(new_n953_), .C2(new_n955_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n445_), .A2(new_n462_), .A3(new_n369_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n913_), .A2(new_n961_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n963_), .A2(G197gat), .A3(new_n762_), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n964_), .A2(KEYINPUT127), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(KEYINPUT127), .ZN(new_n966_));
  AOI21_X1  g765(.A(G197gat), .B1(new_n963_), .B2(new_n762_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n965_), .A2(new_n966_), .A3(new_n967_), .ZN(G1352gat));
  NAND2_X1  g767(.A1(new_n963_), .A2(new_n671_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g769(.A1(new_n963_), .A2(new_n573_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  AND2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n971_), .A2(new_n972_), .A3(new_n973_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n974_), .B1(new_n971_), .B2(new_n972_), .ZN(G1354gat));
  OAI21_X1  g774(.A(G218gat), .B1(new_n962_), .B2(new_n643_), .ZN(new_n976_));
  OR2_X1    g775(.A1(new_n678_), .A2(G218gat), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n962_), .B2(new_n977_), .ZN(G1355gat));
endmodule


