//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT80), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(new_n210_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n205_), .B1(new_n206_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  MUX2_X1   g017(.A(new_n217_), .B(new_n216_), .S(new_n218_), .Z(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(new_n209_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT79), .B1(new_n222_), .B2(G190gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n221_), .B(new_n223_), .C1(new_n224_), .C2(KEYINPUT79), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n215_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G71gat), .B(G99gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G43gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n227_), .B(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G127gat), .B(G134gat), .Z(new_n231_));
  XOR2_X1   g030(.A(G113gat), .B(G120gat), .Z(new_n232_));
  XOR2_X1   g031(.A(new_n231_), .B(new_n232_), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n230_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G227gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(G15gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n234_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT85), .B(G197gat), .ZN(new_n243_));
  INV_X1    g042(.A(G204gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT21), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G211gat), .B(G218gat), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n244_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(G197gat), .B2(G204gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT86), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n248_), .A2(KEYINPUT87), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT21), .B1(new_n248_), .B2(KEYINPUT87), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n245_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT22), .B(G169gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT93), .ZN(new_n261_));
  INV_X1    g060(.A(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n263_), .B(new_n264_), .C1(new_n206_), .C2(new_n209_), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n224_), .B(KEYINPUT92), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n221_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n214_), .A2(new_n219_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT20), .B1(new_n259_), .B2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n215_), .A2(new_n226_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT19), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n271_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT20), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n259_), .B2(new_n270_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n252_), .B(KEYINPUT86), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(new_n257_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n272_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n277_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G8gat), .B(G36gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n265_), .A2(new_n269_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT20), .B1(new_n281_), .B2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n259_), .A2(new_n227_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n293_), .A2(new_n275_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n278_), .B1(new_n281_), .B2(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n259_), .A2(new_n227_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n277_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT32), .B(new_n289_), .C1(new_n295_), .C2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G155gat), .B(G162gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT84), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT3), .Z(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT2), .Z(new_n307_));
  OAI21_X1  g106(.A(new_n303_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n309_));
  AND2_X1   g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(KEYINPUT1), .B2(new_n301_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n233_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n315_), .A2(KEYINPUT4), .ZN(new_n316_));
  INV_X1    g115(.A(new_n233_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n313_), .A3(new_n308_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n318_), .A3(KEYINPUT4), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n300_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G85gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT0), .B(G57gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n300_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n320_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n324_), .B1(new_n320_), .B2(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n291_), .A2(new_n299_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT95), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT33), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n289_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n276_), .B2(new_n283_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n275_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n296_), .A2(new_n277_), .A3(new_n297_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n289_), .A3(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n316_), .A2(new_n300_), .A3(new_n319_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n324_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n315_), .A2(new_n318_), .A3(new_n325_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n338_), .A2(new_n341_), .A3(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n330_), .B1(new_n336_), .B2(new_n346_), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n314_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT28), .B1(new_n314_), .B2(KEYINPUT29), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G22gat), .B(G50gat), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G78gat), .B(G106gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT89), .Z(new_n355_));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n314_), .A2(KEYINPUT29), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n281_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n356_), .B(new_n357_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n259_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n355_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n353_), .B1(new_n364_), .B2(KEYINPUT90), .ZN(new_n365_));
  INV_X1    g164(.A(new_n355_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n363_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n259_), .A2(new_n359_), .B1(new_n357_), .B2(new_n356_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n361_), .A2(new_n355_), .A3(new_n363_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n365_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n370_), .A3(new_n353_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT91), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n369_), .A2(new_n353_), .A3(new_n370_), .A4(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n347_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n329_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n338_), .A2(new_n341_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n289_), .B(KEYINPUT96), .Z(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT27), .A3(new_n341_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n378_), .A2(new_n381_), .A3(new_n384_), .A4(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n241_), .B1(new_n380_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n387_), .ZN(new_n390_));
  NOR4_X1   g189(.A1(new_n390_), .A2(new_n378_), .A3(new_n329_), .A4(new_n240_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G230gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT64), .Z(new_n394_));
  XNOR2_X1  g193(.A(G57gat), .B(G64gat), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n395_), .A2(KEYINPUT11), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(KEYINPUT11), .ZN(new_n397_));
  XOR2_X1   g196(.A(G71gat), .B(G78gat), .Z(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n397_), .A2(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G99gat), .A2(G106gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT6), .ZN(new_n403_));
  OR2_X1    g202(.A1(G85gat), .A2(G92gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G85gat), .A2(G92gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(KEYINPUT9), .A3(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT68), .B(G85gat), .ZN(new_n407_));
  INV_X1    g206(.A(G92gat), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(KEYINPUT9), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n403_), .B(new_n406_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT65), .ZN(new_n412_));
  NAND2_X1  g211(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n412_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT10), .ZN(new_n417_));
  INV_X1    g216(.A(G99gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(KEYINPUT65), .A3(new_n413_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT66), .B(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT67), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n425_));
  AOI211_X1 g224(.A(new_n425_), .B(new_n422_), .C1(new_n416_), .C2(new_n420_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n411_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n404_), .A2(new_n405_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT70), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT8), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n402_), .B(new_n432_), .ZN(new_n433_));
  OR3_X1    g232(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n428_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n403_), .A2(new_n435_), .A3(new_n434_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n439_), .A2(new_n430_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n427_), .A2(KEYINPUT69), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n414_), .A2(new_n415_), .A3(new_n412_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT65), .B1(new_n419_), .B2(new_n413_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n423_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n425_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n421_), .A2(KEYINPUT67), .A3(new_n423_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n410_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n401_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n394_), .B1(new_n450_), .B2(KEYINPUT71), .ZN(new_n451_));
  INV_X1    g250(.A(new_n401_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n438_), .A2(new_n440_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n427_), .A2(KEYINPUT69), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n441_), .A2(new_n401_), .A3(new_n449_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n451_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT12), .B(new_n452_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n394_), .A3(new_n464_), .A4(new_n458_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G120gat), .B(G148gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT5), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G176gat), .B(G204gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n472_));
  INV_X1    g271(.A(new_n470_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n460_), .A2(new_n465_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(KEYINPUT73), .A3(new_n470_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT13), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(KEYINPUT13), .A3(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G8gat), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G29gat), .B(G36gat), .Z(new_n491_));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n490_), .A2(KEYINPUT77), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495_));
  INV_X1    g294(.A(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n488_), .A2(new_n489_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n494_), .A2(new_n498_), .B1(new_n497_), .B2(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n493_), .B(KEYINPUT15), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n497_), .A2(new_n503_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G113gat), .B(G141gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT78), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n502_), .B(new_n511_), .C1(new_n501_), .C2(new_n504_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n481_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n392_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n503_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT34), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n441_), .A2(new_n449_), .A3(new_n493_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n516_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n519_), .A2(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT75), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n516_), .A2(new_n522_), .A3(new_n527_), .A4(new_n521_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n530_));
  XOR2_X1   g329(.A(G190gat), .B(G218gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT74), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n525_), .A2(new_n536_), .A3(new_n528_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n530_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT37), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT37), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n497_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n452_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n490_), .A2(new_n546_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n497_), .B1(G231gat), .B2(G233gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n401_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT76), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G127gat), .B(G155gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT16), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n552_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n548_), .A2(new_n551_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n557_), .B1(new_n560_), .B2(KEYINPUT76), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT17), .B1(new_n560_), .B2(new_n557_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n559_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n545_), .A2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n515_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(new_n483_), .A3(new_n329_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT97), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT38), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n335_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n334_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n338_), .A2(new_n341_), .A3(new_n345_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n284_), .A2(new_n290_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n573_), .A2(new_n574_), .B1(new_n575_), .B2(new_n299_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n388_), .B1(new_n576_), .B2(new_n378_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n240_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n391_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n561_), .A2(new_n562_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n559_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n583_), .A3(new_n540_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n514_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT98), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n587_), .A2(new_n329_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n569_), .B(new_n570_), .C1(new_n483_), .C2(new_n588_), .ZN(G1324gat));
  NAND3_X1  g388(.A1(new_n565_), .A2(new_n484_), .A3(new_n390_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n390_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n584_), .A2(new_n591_), .A3(new_n514_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT99), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n484_), .B1(new_n592_), .B2(KEYINPUT99), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n590_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT40), .B(new_n590_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1325gat));
  AOI21_X1  g401(.A(new_n236_), .B1(new_n587_), .B2(new_n241_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT41), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n565_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(G1326gat));
  INV_X1    g405(.A(G22gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n587_), .B2(new_n378_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n565_), .A2(new_n607_), .A3(new_n378_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1327gat));
  INV_X1    g411(.A(new_n540_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n563_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT103), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n515_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G29gat), .B1(new_n616_), .B2(new_n329_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n580_), .A2(KEYINPUT101), .A3(new_n618_), .A4(new_n545_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n545_), .B(new_n618_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT43), .B1(new_n392_), .B2(new_n544_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n514_), .A2(new_n583_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT102), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT44), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(new_n629_), .A3(new_n625_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n624_), .A2(KEYINPUT44), .A3(new_n625_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n329_), .A2(G29gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n617_), .B1(new_n634_), .B2(new_n635_), .ZN(G1328gat));
  INV_X1    g435(.A(KEYINPUT46), .ZN(new_n637_));
  INV_X1    g436(.A(G36gat), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n390_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n631_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n616_), .A2(new_n638_), .A3(new_n390_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT45), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n637_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT44), .B1(new_n626_), .B2(KEYINPUT102), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n639_), .B1(new_n646_), .B2(new_n630_), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT46), .B(new_n643_), .C1(new_n647_), .C2(new_n638_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(G1329gat));
  NAND2_X1  g448(.A1(new_n241_), .A2(G43gat), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n624_), .A2(KEYINPUT44), .A3(new_n625_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n650_), .B(new_n651_), .C1(new_n646_), .C2(new_n630_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G43gat), .B1(new_n616_), .B2(new_n241_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT47), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT47), .ZN(new_n655_));
  INV_X1    g454(.A(new_n653_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n655_), .B(new_n656_), .C1(new_n633_), .C2(new_n650_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(G1330gat));
  NAND2_X1  g457(.A1(new_n378_), .A2(G50gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n659_), .B(new_n651_), .C1(new_n646_), .C2(new_n630_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G50gat), .B1(new_n616_), .B2(new_n378_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT104), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663_));
  INV_X1    g462(.A(new_n661_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n663_), .B(new_n664_), .C1(new_n633_), .C2(new_n659_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1331gat));
  INV_X1    g465(.A(new_n481_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n513_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n392_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(new_n564_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G57gat), .B1(new_n671_), .B2(new_n329_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n584_), .A2(new_n669_), .ZN(new_n673_));
  INV_X1    g472(.A(G57gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n329_), .B2(KEYINPUT105), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(KEYINPUT105), .B2(new_n674_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n672_), .B1(new_n673_), .B2(new_n676_), .ZN(G1332gat));
  INV_X1    g476(.A(G64gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n673_), .B2(new_n390_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n671_), .A2(new_n678_), .A3(new_n390_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1333gat));
  INV_X1    g482(.A(G71gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n673_), .B2(new_n241_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n671_), .A2(new_n684_), .A3(new_n241_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1334gat));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n673_), .B2(new_n378_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n671_), .A2(new_n690_), .A3(new_n378_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1335gat));
  AND2_X1   g494(.A1(new_n670_), .A2(new_n615_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n329_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n669_), .A2(new_n583_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n624_), .A2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n381_), .A2(new_n407_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(G1336gat));
  NAND3_X1  g500(.A1(new_n696_), .A2(new_n408_), .A3(new_n390_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n699_), .A2(new_n390_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n408_), .ZN(G1337gat));
  NAND3_X1  g503(.A1(new_n696_), .A2(new_n421_), .A3(new_n241_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n699_), .A2(new_n241_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G99gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g510(.A1(new_n696_), .A2(new_n423_), .A3(new_n378_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n624_), .A2(new_n378_), .A3(new_n698_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G106gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G106gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n583_), .B2(new_n668_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n563_), .A2(KEYINPUT110), .A3(new_n513_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n475_), .A2(KEYINPUT13), .A3(new_n476_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT13), .B1(new_n475_), .B2(new_n476_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n722_), .B(KEYINPUT111), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n544_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n481_), .B2(new_n722_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(KEYINPUT112), .A2(KEYINPUT54), .ZN(new_n728_));
  NAND2_X1  g527(.A1(KEYINPUT112), .A2(KEYINPUT54), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n726_), .A2(new_n727_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n734_), .A2(new_n544_), .A3(new_n725_), .A4(new_n729_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n731_), .A2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n464_), .B(new_n458_), .C1(new_n450_), .C2(new_n461_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n394_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n465_), .A2(new_n743_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n454_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n456_), .B2(new_n462_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n746_), .A2(KEYINPUT55), .A3(new_n394_), .A4(new_n464_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n738_), .A2(KEYINPUT113), .A3(new_n739_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n742_), .A2(new_n744_), .A3(new_n747_), .A4(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n470_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(KEYINPUT56), .A3(new_n470_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n509_), .B1(new_n504_), .B2(new_n501_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n499_), .A2(new_n501_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n505_), .A2(new_n509_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n474_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT116), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n474_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n737_), .B1(new_n754_), .B2(new_n762_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n749_), .A2(KEYINPUT56), .A3(new_n470_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT56), .B1(new_n749_), .B2(new_n470_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n737_), .B(new_n762_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n545_), .B1(new_n763_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n475_), .A2(new_n476_), .A3(new_n757_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n475_), .A2(KEYINPUT115), .A3(new_n476_), .A4(new_n757_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n752_), .A2(new_n777_), .A3(new_n753_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n474_), .A2(new_n513_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n764_), .B2(KEYINPUT114), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n776_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n771_), .B1(new_n781_), .B2(new_n613_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n780_), .A2(new_n778_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT57), .B(new_n540_), .C1(new_n783_), .C2(new_n776_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n545_), .B(KEYINPUT118), .C1(new_n763_), .C2(new_n767_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n770_), .A2(new_n782_), .A3(new_n784_), .A4(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n736_), .B1(new_n786_), .B2(new_n563_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n591_), .A2(new_n329_), .A3(new_n379_), .A4(new_n241_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT119), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n513_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT59), .B1(new_n787_), .B2(new_n789_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n782_), .A2(new_n784_), .A3(new_n768_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n563_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n736_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n792_), .A2(KEYINPUT120), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT120), .B1(new_n792_), .B2(new_n798_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n513_), .A2(G113gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n791_), .B1(new_n801_), .B2(new_n802_), .ZN(G1340gat));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n481_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n790_), .B(new_n805_), .C1(KEYINPUT60), .C2(new_n804_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n792_), .A2(new_n667_), .A3(new_n798_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n804_), .ZN(G1341gat));
  AOI21_X1  g607(.A(G127gat), .B1(new_n790_), .B2(new_n583_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n583_), .A2(G127gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n801_), .B2(new_n810_), .ZN(G1342gat));
  AOI21_X1  g610(.A(G134gat), .B1(new_n790_), .B2(new_n613_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n545_), .A2(G134gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n801_), .B2(new_n813_), .ZN(G1343gat));
  NAND2_X1  g613(.A1(new_n786_), .A2(new_n563_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n795_), .ZN(new_n816_));
  NOR4_X1   g615(.A1(new_n379_), .A2(new_n390_), .A3(new_n241_), .A4(new_n381_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n513_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n667_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g621(.A1(new_n816_), .A2(new_n583_), .A3(new_n817_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT121), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n816_), .A2(new_n825_), .A3(new_n583_), .A4(new_n817_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n824_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1346gat));
  AOI21_X1  g629(.A(G162gat), .B1(new_n818_), .B2(new_n613_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n545_), .A2(G162gat), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT122), .Z(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n818_), .B2(new_n833_), .ZN(G1347gat));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n736_), .B1(new_n563_), .B2(new_n793_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n240_), .A2(new_n329_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n379_), .A2(new_n837_), .A3(new_n390_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n836_), .A2(new_n668_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n840_));
  OAI21_X1  g639(.A(G169gat), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n838_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n796_), .A2(new_n513_), .A3(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(KEYINPUT123), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n835_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n204_), .B1(new_n843_), .B2(KEYINPUT123), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(KEYINPUT62), .C1(KEYINPUT123), .C2(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n261_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n847_), .A3(new_n848_), .ZN(G1348gat));
  NOR2_X1   g648(.A1(new_n836_), .A2(new_n838_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G176gat), .B1(new_n850_), .B2(new_n667_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n787_), .A2(new_n838_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(G176gat), .A3(new_n667_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n853_), .A2(KEYINPUT124), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(KEYINPUT124), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n854_), .B2(new_n855_), .ZN(G1349gat));
  AOI21_X1  g655(.A(G183gat), .B1(new_n852_), .B2(new_n583_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n563_), .A2(new_n221_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n850_), .B2(new_n858_), .ZN(G1350gat));
  NAND3_X1  g658(.A1(new_n850_), .A2(new_n613_), .A3(new_n266_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n836_), .A2(new_n544_), .A3(new_n838_), .ZN(new_n861_));
  INV_X1    g660(.A(G190gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(G1351gat));
  NAND3_X1  g662(.A1(new_n378_), .A2(new_n381_), .A3(new_n240_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n390_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n865_), .B2(new_n864_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n816_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n668_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT126), .B(G197gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1352gat));
  NOR2_X1   g670(.A1(new_n868_), .A2(new_n481_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n244_), .A2(KEYINPUT127), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n244_), .A2(KEYINPUT127), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n872_), .B2(new_n874_), .ZN(G1353gat));
  NOR2_X1   g675(.A1(new_n868_), .A2(new_n563_), .ZN(new_n877_));
  OR2_X1    g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT63), .B(G211gat), .Z(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n877_), .B2(new_n880_), .ZN(G1354gat));
  OAI21_X1  g680(.A(G218gat), .B1(new_n868_), .B2(new_n544_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n540_), .A2(G218gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n868_), .B2(new_n883_), .ZN(G1355gat));
endmodule


