//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT82), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n206_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n211_));
  OR2_X1    g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(KEYINPUT22), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT22), .B(G169gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n214_), .B(new_n217_), .C1(new_n218_), .C2(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n213_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT78), .A3(G183gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n227_));
  INV_X1    g026(.A(G183gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT25), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT79), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n224_), .A2(new_n225_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n229_), .A4(new_n223_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT80), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(G169gat), .B2(G176gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n207_), .A2(new_n209_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n237_), .A2(new_n239_), .A3(KEYINPUT24), .A4(new_n220_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n221_), .B1(new_n235_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT30), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G99gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G43gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n249_), .B(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT31), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n253_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n255_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n205_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n259_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n257_), .A3(new_n204_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT0), .ZN(new_n266_));
  INV_X1    g065(.A(G57gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G85gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT96), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G155gat), .ZN(new_n274_));
  INV_X1    g073(.A(G162gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT83), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(G155gat), .B2(G162gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n279_), .B1(new_n283_), .B2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n290_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT2), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT86), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n294_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(KEYINPUT87), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n291_), .A2(KEYINPUT85), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT3), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n291_), .A2(KEYINPUT85), .A3(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n299_), .A2(new_n304_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n278_), .A2(new_n276_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT88), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n293_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n293_), .B2(new_n311_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n204_), .A2(KEYINPUT4), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n273_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n279_), .B1(new_n281_), .B2(new_n280_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n297_), .A2(KEYINPUT86), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n295_), .A2(KEYINPUT2), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n290_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322_));
  NOR4_X1   g121(.A1(new_n322_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n307_), .B1(new_n291_), .B2(KEYINPUT85), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n321_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n318_), .B1(new_n325_), .B2(new_n304_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n292_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n282_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n286_), .A2(KEYINPUT1), .A3(new_n287_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n330_), .B2(new_n279_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT88), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n293_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n205_), .A3(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n289_), .A2(new_n292_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n204_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(KEYINPUT4), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n273_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT97), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT97), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n334_), .A2(new_n340_), .A3(new_n336_), .A4(new_n273_), .ZN(new_n341_));
  AOI221_X4 g140(.A(new_n270_), .B1(new_n317_), .B2(new_n337_), .C1(new_n339_), .C2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n270_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n317_), .A2(new_n337_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT19), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT21), .ZN(new_n351_));
  INV_X1    g150(.A(G211gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(G218gat), .ZN(new_n353_));
  INV_X1    g152(.A(G218gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(G211gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G197gat), .B(G204gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(G211gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(G218gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(KEYINPUT21), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n357_), .A2(KEYINPUT21), .A3(new_n359_), .A4(new_n360_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n362_), .A2(KEYINPUT89), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT89), .B1(new_n362_), .B2(new_n363_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT20), .B1(new_n366_), .B2(new_n246_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n356_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n363_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n241_), .A2(KEYINPUT92), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT24), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n373_), .A3(new_n236_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n210_), .A2(new_n211_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT93), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n210_), .A2(new_n211_), .A3(new_n374_), .A4(KEYINPUT93), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n232_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n371_), .A2(new_n373_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n381_), .A2(new_n220_), .A3(new_n239_), .A4(new_n237_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n243_), .A2(new_n212_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT94), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n218_), .B(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n220_), .B(new_n384_), .C1(new_n386_), .C2(G176gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n370_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n350_), .B1(new_n367_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n362_), .A2(KEYINPUT89), .A3(new_n363_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n246_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n383_), .A2(new_n387_), .A3(new_n370_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .A4(new_n349_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT18), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n349_), .B1(new_n367_), .B2(new_n388_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .A4(new_n350_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n400_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(KEYINPUT27), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT95), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n402_), .A2(new_n407_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  INV_X1    g209(.A(new_n246_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n391_), .A2(new_n392_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n388_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n350_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n403_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n400_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n407_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n409_), .B1(new_n418_), .B2(new_n405_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n347_), .B(new_n406_), .C1(KEYINPUT27), .C2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n332_), .A2(KEYINPUT29), .A3(new_n333_), .ZN(new_n421_));
  AND2_X1   g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n412_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424_));
  OAI22_X1  g223(.A1(new_n335_), .A2(new_n424_), .B1(new_n369_), .B2(new_n368_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n421_), .A2(new_n423_), .B1(new_n425_), .B2(new_n422_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT90), .Z(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT28), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n332_), .A2(new_n333_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n433_), .B2(new_n424_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n432_), .A3(new_n424_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G22gat), .B(G50gat), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n436_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n437_), .B1(new_n440_), .B2(new_n434_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n431_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n428_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n426_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n426_), .B(new_n428_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(new_n431_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n264_), .A2(new_n420_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n344_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n344_), .A2(KEYINPUT33), .A3(new_n343_), .A4(new_n345_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n404_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n405_), .B1(new_n457_), .B2(KEYINPUT95), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n334_), .A2(KEYINPUT4), .A3(new_n336_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n332_), .A2(new_n333_), .A3(new_n316_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n273_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT98), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n337_), .A2(new_n463_), .A3(new_n273_), .A4(new_n460_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n334_), .A2(new_n336_), .A3(new_n272_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n465_), .A2(new_n270_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n467_), .A3(new_n408_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT99), .B1(new_n456_), .B2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n458_), .A2(new_n467_), .A3(new_n408_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT99), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n344_), .A2(new_n345_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n270_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n452_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT101), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n400_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n396_), .B2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n389_), .A2(new_n476_), .A3(new_n395_), .A4(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n402_), .A2(new_n403_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n478_), .B(KEYINPUT100), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n475_), .A2(new_n484_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n469_), .A2(new_n472_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n263_), .B1(new_n420_), .B2(new_n449_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n486_), .A2(new_n487_), .A3(KEYINPUT102), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT102), .B1(new_n486_), .B2(new_n487_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n451_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT6), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  OR3_X1    g292(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G85gat), .B(G92gat), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT8), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT10), .B(G99gat), .Z(new_n499_));
  INV_X1    g298(.A(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G85gat), .A2(G92gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n492_), .B1(KEYINPUT9), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(KEYINPUT9), .B2(new_n496_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n498_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n510_));
  XOR2_X1   g309(.A(G71gat), .B(G78gat), .Z(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n511_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT65), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n508_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n498_), .A2(new_n507_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n515_), .B(KEYINPUT65), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(G230gat), .A3(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n507_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n503_), .A2(new_n506_), .A3(KEYINPUT66), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n498_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n515_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(KEYINPUT12), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n524_), .A2(new_n530_), .A3(new_n531_), .A4(new_n517_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G120gat), .B(G148gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n533_), .A2(new_n537_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT13), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n538_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G169gat), .B(G197gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT73), .B(G8gat), .ZN(new_n551_));
  INV_X1    g350(.A(G1gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n555_), .B(KEYINPUT74), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G29gat), .B(G36gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n563_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n563_), .A2(new_n566_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n566_), .B(KEYINPUT15), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n560_), .A2(new_n562_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n569_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n550_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT77), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n549_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n571_), .A2(new_n576_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT76), .B1(new_n549_), .B2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n546_), .A2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n490_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n518_), .A2(new_n567_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT69), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT35), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n528_), .A2(new_n573_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n592_), .A2(new_n589_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n588_), .A2(new_n597_), .A3(new_n593_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G190gat), .B(G218gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT70), .ZN(new_n600_));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT72), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n598_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n602_), .B(KEYINPUT36), .Z(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n563_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n529_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n515_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n615_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n614_), .A2(new_n516_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n613_), .A2(new_n519_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n620_), .B(KEYINPUT17), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n611_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n585_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n347_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n634_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n596_), .A2(new_n598_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n609_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(KEYINPUT37), .A3(new_n607_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n629_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT75), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n486_), .A2(new_n487_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n486_), .A2(new_n487_), .A3(KEYINPUT102), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n450_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n545_), .B(KEYINPUT67), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR4_X1   g448(.A1(new_n642_), .A2(new_n647_), .A3(new_n583_), .A4(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n552_), .A3(new_n475_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n633_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(KEYINPUT103), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(KEYINPUT103), .ZN(new_n654_));
  OAI221_X1 g453(.A(new_n632_), .B1(new_n633_), .B2(new_n651_), .C1(new_n653_), .C2(new_n654_), .ZN(G1324gat));
  OR2_X1    g454(.A1(new_n419_), .A2(KEYINPUT27), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n406_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n650_), .A2(new_n657_), .A3(new_n551_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n585_), .A2(new_n657_), .A3(new_n630_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G8gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT104), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n663_), .A3(G8gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(KEYINPUT105), .ZN(new_n667_));
  INV_X1    g466(.A(new_n664_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n663_), .B1(new_n659_), .B2(G8gat), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT105), .B(KEYINPUT39), .C1(new_n668_), .C2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n658_), .B1(new_n667_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n673_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n658_), .B(new_n675_), .C1(new_n667_), .C2(new_n671_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n631_), .B2(new_n264_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n650_), .A2(new_n251_), .A3(new_n263_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  OAI21_X1  g481(.A(G22gat), .B1(new_n631_), .B2(new_n448_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  INV_X1    g483(.A(G22gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n650_), .A2(new_n685_), .A3(new_n449_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT107), .Z(G1327gat));
  INV_X1    g487(.A(new_n611_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n628_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n585_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n475_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n608_), .A2(new_n610_), .A3(new_n634_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT37), .B1(new_n638_), .B2(new_n607_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n647_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n490_), .A2(new_n697_), .A3(new_n640_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n584_), .A2(new_n629_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT44), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n703_), .B(new_n700_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n475_), .A2(G29gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n692_), .B1(new_n705_), .B2(new_n706_), .ZN(G1328gat));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n691_), .A2(new_n708_), .A3(new_n657_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT108), .B1(new_n705_), .B2(new_n657_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n490_), .A2(new_n697_), .A3(new_n640_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n697_), .B1(new_n490_), .B2(new_n640_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n701_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n703_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n701_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n716_), .A2(KEYINPUT108), .A3(new_n657_), .A4(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n711_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT110), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(KEYINPUT110), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n716_), .A2(new_n717_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n657_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(G36gat), .A3(new_n718_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n729_), .A2(KEYINPUT110), .A3(new_n721_), .A4(new_n711_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n724_), .A2(new_n730_), .ZN(G1329gat));
  OAI21_X1  g530(.A(G43gat), .B1(new_n726_), .B2(new_n264_), .ZN(new_n732_));
  INV_X1    g531(.A(G43gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n691_), .A2(new_n733_), .A3(new_n263_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n691_), .B2(new_n449_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n449_), .A2(G50gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n705_), .B2(new_n738_), .ZN(G1331gat));
  INV_X1    g538(.A(new_n583_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n642_), .A2(new_n740_), .A3(new_n545_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n490_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n743_), .A2(KEYINPUT111), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(KEYINPUT111), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n475_), .A3(new_n745_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n647_), .A2(new_n740_), .A3(new_n648_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n630_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n347_), .A2(new_n267_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n746_), .A2(new_n267_), .B1(new_n748_), .B2(new_n749_), .ZN(G1332gat));
  INV_X1    g549(.A(G64gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n748_), .B2(new_n657_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n743_), .A2(new_n751_), .A3(new_n657_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1333gat));
  NAND2_X1  g555(.A1(new_n748_), .A2(new_n263_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G71gat), .ZN(new_n758_));
  XOR2_X1   g557(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n759_));
  OR2_X1    g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n742_), .A2(G71gat), .A3(new_n264_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(G1334gat));
  INV_X1    g562(.A(G78gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n748_), .B2(new_n449_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT50), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n743_), .A2(new_n764_), .A3(new_n449_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1335gat));
  AND2_X1   g567(.A1(new_n747_), .A2(new_n690_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n475_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n770_), .A2(KEYINPUT114), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n713_), .A2(new_n714_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n546_), .A2(new_n629_), .A3(new_n583_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(G85gat), .A3(new_n475_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(KEYINPUT114), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n771_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT115), .Z(G1336gat));
  INV_X1    g577(.A(G92gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n769_), .A2(new_n779_), .A3(new_n657_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n772_), .A2(new_n727_), .A3(new_n773_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n779_), .ZN(G1337gat));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n263_), .A2(new_n499_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n769_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n774_), .A2(new_n263_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G99gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G99gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g590(.A1(new_n769_), .A2(new_n500_), .A3(new_n449_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n774_), .A2(new_n449_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G106gat), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT52), .B(new_n500_), .C1(new_n774_), .C2(new_n449_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g597(.A1(new_n657_), .A2(new_n264_), .A3(new_n347_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n575_), .A2(KEYINPUT121), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n575_), .A2(KEYINPUT121), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n569_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n568_), .A2(new_n570_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n549_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n549_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n580_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n542_), .A2(new_n538_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(KEYINPUT122), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n808_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n524_), .A2(new_n530_), .A3(new_n517_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT55), .A3(new_n531_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n532_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n814_), .B(new_n816_), .C1(new_n531_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n537_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT56), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n740_), .A3(new_n542_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n819_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n809_), .B(new_n812_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n689_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT57), .B1(new_n823_), .B2(new_n689_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n818_), .A2(KEYINPUT56), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n817_), .A2(new_n828_), .A3(new_n537_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n827_), .A2(new_n542_), .A3(new_n829_), .A4(new_n807_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n695_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n831_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n640_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT123), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n628_), .B1(new_n826_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n635_), .A2(new_n545_), .A3(new_n639_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n740_), .B2(new_n629_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n583_), .A2(KEYINPUT118), .A3(new_n628_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n841_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n844_), .A2(new_n845_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT119), .B(KEYINPUT54), .C1(new_n849_), .C2(new_n842_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n847_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n448_), .B(new_n799_), .C1(new_n840_), .C2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n853_), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT124), .B1(new_n853_), .B2(KEYINPUT59), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n740_), .B(new_n856_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(G113gat), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n853_), .A2(G113gat), .A3(new_n583_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1340gat));
  OAI211_X1 g661(.A(new_n649_), .B(new_n856_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G120gat), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865_));
  INV_X1    g664(.A(G120gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n546_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n854_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n869_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n853_), .B2(new_n629_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT125), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n874_), .B(new_n871_), .C1(new_n853_), .C2(new_n629_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n858_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n853_), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n877_), .A2(new_n878_), .B1(new_n855_), .B2(new_n854_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n629_), .A2(new_n871_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(G1342gat));
  OAI211_X1 g680(.A(new_n640_), .B(new_n856_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G134gat), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n853_), .A2(G134gat), .A3(new_n689_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1343gat));
  NAND2_X1  g684(.A1(new_n826_), .A2(new_n839_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n852_), .B1(new_n886_), .B2(new_n629_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n263_), .A2(new_n448_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n887_), .A2(new_n347_), .A3(new_n657_), .A4(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n740_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n649_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n890_), .A2(new_n628_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  NAND3_X1  g696(.A1(new_n890_), .A2(new_n275_), .A3(new_n611_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n890_), .A2(new_n640_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n275_), .ZN(G1347gat));
  INV_X1    g699(.A(new_n887_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n727_), .A2(new_n475_), .A3(new_n264_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n448_), .A3(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903_), .B2(new_n583_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(G169gat), .C1(new_n903_), .C2(new_n583_), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n903_), .A2(new_n386_), .A3(new_n583_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1348gat));
  OAI21_X1  g708(.A(G176gat), .B1(new_n903_), .B2(new_n648_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n546_), .A2(new_n214_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n903_), .B2(new_n911_), .ZN(G1349gat));
  NOR2_X1   g711(.A1(new_n903_), .A2(new_n629_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n379_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n228_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n903_), .B2(new_n695_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n611_), .A2(new_n232_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n903_), .B2(new_n917_), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n889_), .A2(new_n727_), .A3(new_n475_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n901_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n583_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT126), .B(G197gat), .Z(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1352gat));
  INV_X1    g722(.A(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n649_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n628_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT63), .B(G211gat), .Z(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1354gat));
  NOR3_X1   g729(.A1(new_n920_), .A2(new_n354_), .A3(new_n695_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n920_), .A2(KEYINPUT127), .A3(new_n689_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(G218gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT127), .B1(new_n920_), .B2(new_n689_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n931_), .B1(new_n933_), .B2(new_n934_), .ZN(G1355gat));
endmodule


