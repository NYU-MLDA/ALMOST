//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_, new_n970_, new_n971_,
    new_n973_, new_n974_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_, new_n990_;
  AND2_X1   g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n207_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT10), .B(G99gat), .Z(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n205_), .A2(new_n219_), .A3(KEYINPUT9), .ZN(new_n220_));
  INV_X1    g019(.A(new_n206_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(new_n219_), .C2(KEYINPUT9), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n205_), .A2(new_n219_), .A3(KEYINPUT9), .A4(new_n206_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n218_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G57gat), .B(G64gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n226_));
  XOR2_X1   g025(.A(G71gat), .B(G78gat), .Z(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n227_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n215_), .A2(new_n224_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT65), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n215_), .A2(new_n224_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n202_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n234_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n202_), .B1(new_n239_), .B2(new_n231_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n236_), .A2(KEYINPUT12), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT12), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n240_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G120gat), .B(G148gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT5), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G176gat), .B(G204gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n238_), .A2(new_n244_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT13), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT66), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(KEYINPUT66), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT105), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(KEYINPUT3), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(KEYINPUT3), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT83), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT83), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(G141gat), .A3(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT2), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT87), .B1(new_n271_), .B2(KEYINPUT86), .ZN(new_n272_));
  INV_X1    g071(.A(new_n263_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n264_), .A2(new_n270_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n282_), .A2(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT85), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT1), .B1(new_n277_), .B2(new_n278_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n285_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n273_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n284_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT98), .ZN(new_n304_));
  INV_X1    g103(.A(new_n300_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n297_), .A2(new_n298_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n299_), .A2(KEYINPUT98), .A3(new_n300_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n307_), .A2(new_n284_), .A3(new_n295_), .A4(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n303_), .A2(KEYINPUT4), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT99), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n301_), .B1(new_n284_), .B2(new_n295_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n303_), .A2(new_n309_), .A3(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G57gat), .B(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n310_), .A2(new_n316_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT104), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n318_), .A2(new_n324_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n318_), .A2(new_n324_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT104), .B1(new_n331_), .B2(new_n317_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n326_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(G183gat), .ZN(new_n338_));
  INV_X1    g137(.A(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G169gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT22), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT22), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n347_), .A2(KEYINPUT96), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT96), .B1(new_n347_), .B2(new_n348_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n341_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT25), .B(G183gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n334_), .A2(KEYINPUT23), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n342_), .A2(new_n346_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(KEYINPUT24), .A3(new_n348_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT24), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n354_), .A2(new_n357_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT95), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n348_), .A2(KEYINPUT24), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n362_), .B1(new_n365_), .B2(new_n360_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n357_), .A4(new_n354_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n351_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(G197gat), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n374_));
  INV_X1    g173(.A(G197gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(G204gat), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT21), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n373_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n373_), .A2(new_n378_), .A3(KEYINPUT92), .A4(new_n381_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n380_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n376_), .A2(new_n377_), .ZN(new_n391_));
  INV_X1    g190(.A(G204gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT91), .B(G204gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n375_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n390_), .B1(new_n396_), .B2(KEYINPUT21), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n384_), .B1(new_n389_), .B2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n370_), .A2(KEYINPUT97), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT97), .B1(new_n370_), .B2(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT19), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n341_), .A2(new_n348_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n347_), .A2(KEYINPUT80), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT22), .B(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n346_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n405_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT25), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT25), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n339_), .A2(KEYINPUT26), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT26), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G190gat), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n412_), .A2(new_n414_), .A3(new_n415_), .A4(new_n417_), .ZN(new_n418_));
  AND4_X1   g217(.A1(new_n418_), .A2(new_n357_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n410_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n404_), .B1(new_n398_), .B2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n399_), .A2(new_n400_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n402_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n389_), .A2(new_n397_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n383_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n351_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n403_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n398_), .A2(new_n420_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n423_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n422_), .A2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G8gat), .B(G36gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT18), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n333_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT103), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n398_), .B2(new_n420_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n413_), .A2(G183gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n338_), .A2(KEYINPUT25), .ZN(new_n442_));
  AND4_X1   g241(.A1(new_n415_), .A2(new_n417_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n355_), .A2(new_n356_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n443_), .A2(new_n366_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n347_), .A2(new_n348_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT96), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n347_), .A2(KEYINPUT96), .A3(new_n348_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n445_), .B1(new_n450_), .B2(new_n341_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n451_), .A2(new_n424_), .A3(new_n383_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n402_), .B1(new_n440_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n425_), .A2(new_n426_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n454_), .A2(KEYINPUT20), .A3(new_n423_), .A4(new_n428_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n435_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n438_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AOI211_X1 g257(.A(KEYINPUT103), .B(new_n435_), .C1(new_n453_), .C2(new_n455_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n258_), .B1(new_n437_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n435_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(new_n438_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n328_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n331_), .A2(KEYINPUT104), .A3(new_n317_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n466_), .A2(new_n326_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n467_), .A3(KEYINPUT105), .ZN(new_n468_));
  INV_X1    g267(.A(new_n434_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT20), .B1(new_n370_), .B2(new_n398_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n428_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n402_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT97), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n398_), .A2(new_n420_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n370_), .A2(KEYINPUT97), .A3(new_n398_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .A4(new_n404_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n473_), .A2(new_n478_), .A3(new_n434_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n303_), .A2(KEYINPUT101), .A3(new_n309_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT101), .B1(new_n303_), .B2(new_n309_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n312_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n312_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n324_), .B1(new_n310_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n331_), .A2(KEYINPUT33), .A3(new_n317_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n480_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n461_), .A2(new_n468_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G228gat), .ZN(new_n494_));
  INV_X1    g293(.A(G233gat), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n495_), .A2(KEYINPUT89), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(KEYINPUT89), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT93), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G22gat), .B(G50gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n504_));
  NOR3_X1   g303(.A1(new_n296_), .A2(KEYINPUT29), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n276_), .A2(new_n283_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n296_), .B2(KEYINPUT29), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n508_), .A3(new_n506_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n502_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n508_), .B1(new_n284_), .B2(new_n295_), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n398_), .A2(new_n515_), .B1(new_n499_), .B2(new_n498_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(G78gat), .ZN(new_n517_));
  INV_X1    g316(.A(G78gat), .ZN(new_n518_));
  OAI221_X1 g317(.A(new_n518_), .B1(new_n499_), .B2(new_n498_), .C1(new_n398_), .C2(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n514_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT94), .B(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(new_n513_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n522_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n493_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n524_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n522_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n521_), .A2(new_n524_), .A3(new_n522_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n333_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n422_), .A2(new_n429_), .A3(new_n469_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT27), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n456_), .A2(new_n469_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT106), .B1(new_n480_), .B2(new_n535_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT106), .ZN(new_n540_));
  AOI211_X1 g339(.A(new_n540_), .B(KEYINPUT27), .C1(new_n470_), .C2(new_n479_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n533_), .B(new_n538_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n528_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(G15gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n348_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n548_));
  NOR2_X1   g347(.A1(G183gat), .A2(G190gat), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n550_), .B2(new_n337_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n408_), .B1(new_n407_), .B2(new_n346_), .ZN(new_n552_));
  AND4_X1   g351(.A1(new_n408_), .A2(new_n343_), .A3(new_n345_), .A4(new_n346_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n418_), .A2(new_n357_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n554_), .A2(KEYINPUT30), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT30), .B1(new_n554_), .B2(new_n555_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G71gat), .B(G99gat), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n410_), .B2(new_n419_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n554_), .A2(KEYINPUT30), .A3(new_n555_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n546_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT81), .B(G43gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n558_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n546_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n565_), .A2(new_n566_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT82), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n566_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT31), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n565_), .A2(new_n570_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n566_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(new_n572_), .A3(new_n571_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n301_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n575_), .A2(new_n302_), .A3(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n575_), .A2(new_n302_), .A3(new_n580_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n302_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n585_), .A2(new_n586_), .A3(new_n333_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n434_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n535_), .B1(new_n534_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n540_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n480_), .A2(KEYINPUT106), .A3(new_n535_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n590_), .A2(new_n591_), .B1(new_n537_), .B2(new_n536_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n587_), .A2(KEYINPUT107), .A3(new_n527_), .A4(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT107), .ZN(new_n594_));
  INV_X1    g393(.A(new_n333_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n582_), .A2(new_n595_), .A3(new_n583_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n527_), .B(new_n538_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n594_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n543_), .A2(new_n584_), .B1(new_n593_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G29gat), .B(G36gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G43gat), .B(G50gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT70), .B(G1gat), .Z(new_n605_));
  INV_X1    g404(.A(G8gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT14), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G15gat), .B(G22gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G1gat), .B(G8gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n604_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT76), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n619_), .A2(new_n620_), .B1(new_n614_), .B2(new_n604_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n604_), .A2(new_n614_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n618_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n621_), .A2(new_n624_), .A3(G229gat), .A4(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n602_), .B(KEYINPUT15), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n613_), .A3(new_n612_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n615_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G113gat), .B(G141gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT77), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT78), .Z(new_n632_));
  XNOR2_X1  g431(.A(G169gat), .B(G197gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n625_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n625_), .B2(new_n629_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n257_), .A2(new_n599_), .A3(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n639_));
  NAND2_X1  g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n234_), .A2(new_n626_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT68), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n239_), .A2(new_n602_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n643_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G190gat), .B(G218gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n646_), .A2(new_n648_), .B1(KEYINPUT36), .B2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n643_), .B(new_n647_), .C1(new_n645_), .C2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n651_), .A2(KEYINPUT36), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n652_), .B(new_n654_), .C1(KEYINPUT36), .C2(new_n651_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(KEYINPUT69), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT37), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n231_), .B(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(new_n614_), .Z(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT71), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n663_), .B(new_n614_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT71), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(G127gat), .B(G155gat), .Z(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT16), .ZN(new_n670_));
  XNOR2_X1  g469(.A(G183gat), .B(G211gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT17), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n665_), .A2(new_n668_), .A3(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT72), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n672_), .A2(new_n673_), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n666_), .A2(new_n674_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT73), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT73), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(new_n681_), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n661_), .A2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n638_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n333_), .A2(new_n605_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT108), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT108), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT38), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n257_), .A2(new_n679_), .A3(new_n637_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n657_), .A2(new_n658_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n599_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G1gat), .B1(new_n698_), .B2(new_n595_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n688_), .A2(KEYINPUT38), .A3(new_n689_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n692_), .A2(new_n699_), .A3(new_n700_), .ZN(G1324gat));
  INV_X1    g500(.A(new_n592_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n685_), .A2(new_n606_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT39), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n697_), .A2(new_n702_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G8gat), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT39), .B(new_n606_), .C1(new_n697_), .C2(new_n702_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT40), .B(new_n703_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1325gat));
  INV_X1    g511(.A(new_n584_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n685_), .A2(new_n545_), .A3(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT109), .Z(new_n715_));
  OAI21_X1  g514(.A(G15gat), .B1(new_n698_), .B2(new_n584_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT41), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n716_), .A2(KEYINPUT41), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n717_), .A3(new_n718_), .ZN(G1326gat));
  INV_X1    g518(.A(G22gat), .ZN(new_n720_));
  INV_X1    g519(.A(new_n527_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n697_), .B2(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT42), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n685_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1327gat));
  INV_X1    g524(.A(new_n683_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n694_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n638_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G29gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n333_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n637_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n255_), .A2(new_n683_), .A3(new_n731_), .A4(new_n256_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n593_), .A2(new_n598_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n333_), .B(new_n436_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n491_), .B1(new_n736_), .B2(new_n258_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n721_), .B1(new_n737_), .B2(new_n468_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n542_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n584_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n735_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n734_), .B1(new_n741_), .B2(new_n661_), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT43), .B(new_n660_), .C1(new_n735_), .C2(new_n740_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n733_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT110), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n599_), .B2(new_n660_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(new_n734_), .A3(new_n661_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n732_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(KEYINPUT44), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n333_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755_));
  OAI21_X1  g554(.A(G29gat), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT44), .B1(new_n744_), .B2(KEYINPUT110), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n757_), .A2(new_n750_), .B1(KEYINPUT44), .B2(new_n748_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT111), .B1(new_n758_), .B2(new_n333_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n730_), .B1(new_n756_), .B2(new_n759_), .ZN(G1328gat));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT114), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT115), .Z(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n257_), .A2(new_n637_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n592_), .A2(G36gat), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(new_n727_), .A3(new_n741_), .A4(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT113), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n767_), .B(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n592_), .B1(new_n748_), .B2(KEYINPUT44), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n751_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT110), .B(new_n732_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n770_), .B1(new_n774_), .B2(G36gat), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n761_), .A2(KEYINPUT114), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n764_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n776_), .ZN(new_n778_));
  INV_X1    g577(.A(G36gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n752_), .B2(new_n771_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n778_), .B(new_n763_), .C1(new_n780_), .C2(new_n770_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n781_), .ZN(G1329gat));
  NAND4_X1  g581(.A1(new_n752_), .A2(G43gat), .A3(new_n713_), .A4(new_n753_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n728_), .A2(new_n713_), .ZN(new_n784_));
  INV_X1    g583(.A(G43gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n783_), .A2(KEYINPUT47), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT47), .B1(new_n783_), .B2(new_n786_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1330gat));
  AOI21_X1  g588(.A(G50gat), .B1(new_n728_), .B2(new_n721_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n721_), .A2(G50gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n758_), .B2(new_n791_), .ZN(G1331gat));
  AND3_X1   g591(.A1(new_n680_), .A2(new_n682_), .A3(new_n637_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n257_), .A2(new_n741_), .A3(new_n694_), .A4(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n333_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n599_), .A2(new_n731_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n798_), .A2(new_n684_), .A3(new_n257_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n595_), .A2(G57gat), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n797_), .A2(G57gat), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT117), .ZN(G1332gat));
  INV_X1    g601(.A(G64gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n796_), .B2(new_n702_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT48), .Z(new_n805_));
  NAND3_X1  g604(.A1(new_n799_), .A2(new_n803_), .A3(new_n702_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1333gat));
  INV_X1    g606(.A(G71gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n796_), .B2(new_n713_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT49), .Z(new_n810_));
  NAND3_X1  g609(.A1(new_n799_), .A2(new_n808_), .A3(new_n713_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1334gat));
  NAND3_X1  g611(.A1(new_n799_), .A2(new_n518_), .A3(new_n721_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n794_), .A2(KEYINPUT116), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n794_), .A2(KEYINPUT116), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n721_), .A3(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(G78gat), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(G78gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT119), .B(new_n813_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1335gat));
  INV_X1    g623(.A(new_n257_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n825_), .A2(new_n726_), .A3(new_n731_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n746_), .A2(new_n747_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G85gat), .B1(new_n829_), .B2(new_n595_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n798_), .A2(new_n257_), .A3(new_n727_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n203_), .A3(new_n333_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1336gat));
  OAI21_X1  g632(.A(G92gat), .B1(new_n829_), .B2(new_n592_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n204_), .A3(new_n702_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1337gat));
  NAND2_X1  g635(.A1(new_n828_), .A2(new_n713_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n713_), .A2(new_n217_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n837_), .A2(G99gat), .B1(new_n831_), .B2(new_n838_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g639(.A1(new_n831_), .A2(new_n216_), .A3(new_n721_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n826_), .A2(new_n827_), .A3(new_n721_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n842_), .A2(new_n843_), .A3(G106gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n842_), .B2(G106gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g646(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n793_), .A2(new_n660_), .A3(new_n254_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n660_), .A2(new_n254_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n680_), .A2(new_n682_), .A3(new_n637_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n253_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n625_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n621_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n628_), .B1(new_n604_), .B2(new_n614_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n634_), .B1(new_n858_), .B2(new_n627_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT121), .B1(new_n855_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n856_), .A2(new_n860_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n253_), .A3(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n241_), .A2(new_n243_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n202_), .B1(new_n866_), .B2(new_n233_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n244_), .A2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(KEYINPUT55), .B(new_n240_), .C1(new_n241_), .C2(new_n243_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n867_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n249_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(KEYINPUT56), .A3(new_n249_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n252_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n862_), .B(new_n865_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n694_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n863_), .A2(new_n252_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n871_), .B2(new_n249_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(KEYINPUT122), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n875_), .B1(new_n883_), .B2(KEYINPUT122), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n882_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n882_), .B(KEYINPUT58), .C1(new_n884_), .C2(new_n885_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n661_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n862_), .A2(new_n865_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n877_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT57), .B(new_n694_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n881_), .A2(new_n890_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n854_), .B1(new_n894_), .B2(new_n683_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n713_), .A2(new_n333_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n597_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n895_), .A2(KEYINPUT59), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n854_), .B1(new_n894_), .B2(new_n679_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT59), .B1(new_n900_), .B2(new_n898_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G113gat), .B1(new_n902_), .B2(new_n637_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n900_), .A2(new_n904_), .A3(new_n898_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n900_), .B2(new_n898_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n637_), .A2(G113gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n903_), .B1(new_n907_), .B2(new_n908_), .ZN(G1340gat));
  OAI21_X1  g708(.A(G120gat), .B1(new_n902_), .B2(new_n825_), .ZN(new_n910_));
  INV_X1    g709(.A(G120gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n825_), .B2(KEYINPUT60), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(KEYINPUT60), .B2(new_n911_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n910_), .B1(new_n907_), .B2(new_n913_), .ZN(G1341gat));
  OAI21_X1  g713(.A(G127gat), .B1(new_n902_), .B2(new_n679_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n683_), .A2(G127gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n907_), .B2(new_n916_), .ZN(G1342gat));
  INV_X1    g716(.A(new_n902_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n661_), .A2(G134gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT124), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n905_), .A2(new_n695_), .A3(new_n906_), .ZN(new_n921_));
  INV_X1    g720(.A(G134gat), .ZN(new_n922_));
  AOI22_X1  g721(.A1(new_n918_), .A2(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1343gat));
  NAND4_X1  g722(.A1(new_n592_), .A2(new_n584_), .A3(new_n333_), .A4(new_n721_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT125), .B1(new_n900_), .B2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n900_), .A2(KEYINPUT125), .A3(new_n924_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G141gat), .B1(new_n928_), .B2(new_n637_), .ZN(new_n929_));
  INV_X1    g728(.A(G141gat), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n930_), .B(new_n731_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1344gat));
  OAI21_X1  g731(.A(G148gat), .B1(new_n928_), .B2(new_n825_), .ZN(new_n933_));
  INV_X1    g732(.A(G148gat), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n934_), .B(new_n257_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1345gat));
  XNOR2_X1  g735(.A(KEYINPUT61), .B(G155gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n928_), .B2(new_n683_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n937_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n726_), .B(new_n939_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1346gat));
  INV_X1    g740(.A(new_n927_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n660_), .B1(new_n942_), .B2(new_n925_), .ZN(new_n943_));
  INV_X1    g742(.A(G162gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n695_), .A2(new_n944_), .ZN(new_n945_));
  OAI22_X1  g744(.A1(new_n943_), .A2(new_n944_), .B1(new_n928_), .B2(new_n945_), .ZN(G1347gat));
  NOR2_X1   g745(.A1(new_n596_), .A2(new_n592_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n721_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n893_), .ZN(new_n950_));
  AOI21_X1  g749(.A(KEYINPUT57), .B1(new_n878_), .B2(new_n694_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n726_), .B1(new_n952_), .B2(new_n890_), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n731_), .B(new_n949_), .C1(new_n953_), .C2(new_n854_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n954_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n955_));
  INV_X1    g754(.A(new_n949_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n895_), .A2(new_n956_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n957_), .A2(new_n407_), .A3(new_n731_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n955_), .A2(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(KEYINPUT62), .B1(new_n954_), .B2(G169gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(KEYINPUT126), .B1(new_n959_), .B2(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n960_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n962_), .A2(new_n963_), .A3(new_n958_), .A4(new_n955_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n961_), .A2(new_n964_), .ZN(G1348gat));
  AOI21_X1  g764(.A(G176gat), .B1(new_n957_), .B2(new_n257_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n900_), .A2(new_n721_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n825_), .A2(new_n346_), .A3(new_n948_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(G1349gat));
  NAND3_X1  g768(.A1(new_n967_), .A2(new_n726_), .A3(new_n947_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n679_), .A2(new_n353_), .ZN(new_n971_));
  AOI22_X1  g770(.A1(new_n970_), .A2(new_n338_), .B1(new_n957_), .B2(new_n971_), .ZN(G1350gat));
  NAND3_X1  g771(.A1(new_n957_), .A2(new_n695_), .A3(new_n352_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n895_), .A2(new_n660_), .A3(new_n956_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n339_), .B2(new_n974_), .ZN(G1351gat));
  NAND3_X1  g774(.A1(new_n702_), .A2(new_n533_), .A3(new_n584_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n900_), .A2(new_n976_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n977_), .A2(new_n731_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g778(.A1(new_n900_), .A2(new_n825_), .A3(new_n976_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n980_), .A2(G204gat), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n394_), .B2(new_n980_), .ZN(G1353gat));
  NAND3_X1  g781(.A1(new_n977_), .A2(new_n676_), .A3(new_n678_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n984_));
  AND2_X1   g783(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n985_));
  NOR3_X1   g784(.A1(new_n983_), .A2(new_n984_), .A3(new_n985_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n986_), .B1(new_n983_), .B2(new_n984_), .ZN(G1354gat));
  INV_X1    g786(.A(G218gat), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n977_), .A2(new_n988_), .A3(new_n695_), .ZN(new_n989_));
  NOR3_X1   g788(.A1(new_n900_), .A2(new_n660_), .A3(new_n976_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n990_), .B2(new_n988_), .ZN(G1355gat));
endmodule


