//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n594_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n208_));
  INV_X1    g007(.A(G197gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT89), .B1(new_n207_), .B2(G197gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT21), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G218gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G211gat), .ZN(new_n215_));
  INV_X1    g014(.A(G211gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G218gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT90), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n209_), .B2(G204gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n207_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n209_), .B2(G204gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n207_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n220_), .B(new_n221_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n213_), .B(new_n218_), .C1(new_n225_), .C2(KEYINPUT21), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT21), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n225_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n227_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n226_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT23), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(KEYINPUT24), .A3(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT26), .B(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n240_), .A2(new_n241_), .B1(new_n242_), .B2(new_n235_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n234_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n237_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n244_), .A2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n232_), .A2(KEYINPUT93), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT22), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(G169gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n249_), .B(new_n256_), .C1(new_n248_), .C2(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n246_), .A2(new_n257_), .A3(new_n237_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n244_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT20), .B1(new_n232_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT93), .B1(new_n232_), .B2(new_n252_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n253_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT19), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n232_), .A2(new_n259_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT20), .B1(new_n232_), .B2(new_n252_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n206_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT101), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n264_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT91), .B1(new_n207_), .B2(G197gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n222_), .A2(new_n209_), .A3(G204gat), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n220_), .A2(new_n221_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n229_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT92), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n225_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(new_n244_), .A3(new_n258_), .A4(new_n226_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n239_), .A2(new_n243_), .B1(new_n246_), .B2(new_n250_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n280_), .B2(new_n226_), .ZN(new_n283_));
  OAI211_X1 g082(.A(KEYINPUT20), .B(new_n281_), .C1(new_n283_), .C2(KEYINPUT93), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n264_), .B1(new_n284_), .B2(new_n253_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT94), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n272_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(KEYINPUT94), .B(new_n264_), .C1(new_n284_), .C2(new_n253_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n206_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n271_), .A2(KEYINPUT27), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT27), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n286_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n272_), .ZN(new_n293_));
  AND4_X1   g092(.A1(new_n206_), .A2(new_n292_), .A3(new_n288_), .A4(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n206_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n291_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G228gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G78gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G106gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G22gat), .B(G50gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  INV_X1    g103(.A(G155gat), .ZN(new_n305_));
  INV_X1    g104(.A(G162gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n308_), .B2(new_n307_), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(KEYINPUT2), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(KEYINPUT3), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT87), .B(KEYINPUT2), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT88), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n313_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n323_), .B2(new_n313_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n322_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n307_), .A2(new_n304_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n317_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n331_), .A2(KEYINPUT28), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n232_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(KEYINPUT28), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n303_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n336_), .A3(new_n302_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT86), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G120gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n345_), .B(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n330_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n330_), .A2(new_n348_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(KEYINPUT4), .A3(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(KEYINPUT4), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(G225gat), .A4(G233gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n349_), .A2(new_n354_), .A3(new_n350_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT97), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n349_), .A2(KEYINPUT97), .A3(new_n354_), .A4(new_n350_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT100), .ZN(new_n365_));
  INV_X1    g164(.A(new_n363_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n353_), .A2(new_n366_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT100), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n359_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G43gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT30), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(new_n259_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT85), .B(G15gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n348_), .B(KEYINPUT31), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n380_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n370_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n297_), .A2(new_n343_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AND4_X1   g185(.A1(KEYINPUT32), .A2(new_n266_), .A3(new_n206_), .A4(new_n269_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n292_), .A2(new_n288_), .A3(new_n293_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(KEYINPUT99), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT99), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n370_), .A2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n349_), .A2(new_n350_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n363_), .B1(new_n396_), .B2(new_n354_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT33), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n367_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n357_), .A2(new_n358_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(KEYINPUT33), .A3(new_n366_), .A4(new_n353_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT96), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n206_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n388_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(KEYINPUT96), .A3(new_n289_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n402_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n394_), .B1(new_n408_), .B2(KEYINPUT98), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n410_));
  AOI211_X1 g209(.A(new_n410_), .B(new_n402_), .C1(new_n404_), .C2(new_n407_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n343_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n370_), .A2(new_n343_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n413_), .A2(new_n296_), .A3(new_n290_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n386_), .B1(new_n416_), .B2(new_n383_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT78), .B(G15gat), .ZN(new_n418_));
  INV_X1    g217(.A(G22gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G1gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G1gat), .B(G8gat), .Z(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n424_), .B(KEYINPUT79), .ZN(new_n429_));
  INV_X1    g228(.A(new_n427_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G29gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT74), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G43gat), .B(G50gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT75), .B(KEYINPUT15), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n436_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G229gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT82), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n432_), .A2(new_n436_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n438_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n446_), .B2(new_n442_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G113gat), .B(G141gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT83), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G169gat), .B(G197gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n451_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n444_), .B(new_n453_), .C1(new_n446_), .C2(new_n442_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n417_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G85gat), .A3(G92gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G85gat), .B(G92gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n465_), .B(KEYINPUT6), .Z(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT10), .B(G99gat), .Z(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT64), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n471_), .A3(new_n468_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n466_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT70), .ZN(new_n475_));
  INV_X1    g274(.A(new_n460_), .ZN(new_n476_));
  OR3_X1    g275(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n476_), .B1(new_n466_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT8), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n440_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT76), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT76), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n485_), .A3(new_n440_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n481_), .B2(new_n474_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n487_), .A3(new_n474_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n436_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n484_), .A2(new_n486_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT34), .Z(new_n496_));
  XNOR2_X1  g295(.A(G190gat), .B(G218gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G134gat), .B(G162gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n494_), .A2(new_n496_), .B1(KEYINPUT36), .B2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n496_), .B(KEYINPUT73), .Z(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT35), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n494_), .B2(KEYINPUT77), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n483_), .A2(KEYINPUT76), .B1(new_n491_), .B2(new_n492_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n486_), .A4(new_n502_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n500_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n499_), .A2(KEYINPUT36), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n500_), .A2(new_n504_), .A3(new_n511_), .A4(new_n507_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT37), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G231gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n432_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G71gat), .B(G78gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(KEYINPUT11), .B2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n519_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n516_), .B(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G127gat), .B(G155gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT16), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G183gat), .B(G211gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n529_), .A2(KEYINPUT80), .A3(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n529_), .A2(new_n530_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n525_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n525_), .A2(new_n531_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT81), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n514_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G230gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n489_), .A2(new_n524_), .A3(new_n490_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n490_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n523_), .B1(new_n543_), .B2(new_n488_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n539_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(KEYINPUT69), .B(new_n539_), .C1(new_n542_), .C2(new_n545_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n540_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n524_), .A2(KEYINPUT12), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n482_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n551_), .A2(new_n554_), .A3(new_n538_), .A4(new_n544_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n548_), .A2(new_n549_), .A3(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G120gat), .B(G148gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT71), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n556_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n537_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n457_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n370_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n569_), .A2(G1gat), .A3(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n571_), .A2(KEYINPUT38), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(KEYINPUT38), .ZN(new_n573_));
  INV_X1    g372(.A(new_n513_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n417_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n567_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n455_), .A3(new_n576_), .A4(new_n535_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G1gat), .B1(new_n577_), .B2(new_n570_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n573_), .A3(new_n578_), .ZN(G1324gat));
  OAI21_X1  g378(.A(G8gat), .B1(new_n577_), .B2(new_n297_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT102), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT102), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT39), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n569_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n297_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n422_), .A3(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n583_), .B(new_n586_), .C1(KEYINPUT39), .C2(new_n582_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT40), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(G1325gat));
  OAI21_X1  g388(.A(G15gat), .B1(new_n577_), .B2(new_n383_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT41), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n569_), .A2(G15gat), .A3(new_n383_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(G1326gat));
  OAI21_X1  g392(.A(G22gat), .B1(new_n577_), .B2(new_n343_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT42), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n584_), .A2(new_n419_), .A3(new_n342_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1327gat));
  INV_X1    g396(.A(new_n536_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n574_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n567_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n457_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(G29gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n370_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT104), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT43), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n513_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n383_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n606_), .B(new_n608_), .C1(new_n610_), .C2(new_n386_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT103), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT43), .B1(new_n417_), .B2(new_n514_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n402_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n406_), .A2(KEYINPUT96), .A3(new_n289_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT96), .B1(new_n406_), .B2(new_n289_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n410_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n408_), .A2(KEYINPUT98), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n394_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n414_), .B1(new_n620_), .B2(new_n343_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n385_), .B1(new_n621_), .B2(new_n609_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n606_), .A4(new_n608_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n612_), .A2(new_n613_), .A3(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n567_), .A2(new_n456_), .A3(new_n536_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT44), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n570_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(KEYINPUT44), .A3(new_n626_), .ZN(new_n630_));
  AOI211_X1 g429(.A(new_n605_), .B(new_n603_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n628_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n370_), .A3(new_n630_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT104), .B1(new_n633_), .B2(G29gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n604_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT105), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n637_), .B(new_n604_), .C1(new_n631_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(G1328gat));
  INV_X1    g438(.A(G36gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n602_), .A2(new_n640_), .A3(new_n585_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT45), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n297_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n644_));
  AOI211_X1 g443(.A(new_n643_), .B(new_n640_), .C1(new_n644_), .C2(new_n630_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n632_), .A2(new_n585_), .A3(new_n630_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT106), .B1(new_n646_), .B2(G36gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT46), .B(new_n642_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  AOI21_X1  g451(.A(G43gat), .B1(new_n602_), .B2(new_n609_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n632_), .A2(G43gat), .A3(new_n609_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n630_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT47), .Z(G1330gat));
  OR3_X1    g455(.A1(new_n601_), .A2(G50gat), .A3(new_n343_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n632_), .A2(new_n342_), .A3(new_n630_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G50gat), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n658_), .A2(new_n659_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(G1331gat));
  NAND4_X1  g462(.A1(new_n575_), .A2(new_n456_), .A3(new_n567_), .A4(new_n536_), .ZN(new_n664_));
  INV_X1    g463(.A(G57gat), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n570_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n417_), .A2(new_n455_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(new_n567_), .A3(new_n536_), .A4(new_n514_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n570_), .B1(new_n668_), .B2(KEYINPUT108), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(KEYINPUT108), .B2(new_n668_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n666_), .B1(new_n670_), .B2(new_n665_), .ZN(G1332gat));
  OAI21_X1  g470(.A(G64gat), .B1(new_n664_), .B2(new_n297_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT48), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n297_), .A2(G64gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n668_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT109), .Z(G1333gat));
  OAI21_X1  g475(.A(G71gat), .B1(new_n664_), .B2(new_n383_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n383_), .A2(G71gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n668_), .B2(new_n680_), .ZN(G1334gat));
  OAI21_X1  g480(.A(G78gat), .B1(new_n664_), .B2(new_n343_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT50), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n343_), .A2(G78gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n668_), .B2(new_n684_), .ZN(G1335gat));
  INV_X1    g484(.A(G85gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n599_), .A2(new_n576_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n667_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(new_n570_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT111), .Z(new_n690_));
  NOR3_X1   g489(.A1(new_n576_), .A2(new_n455_), .A3(new_n536_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n625_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n686_), .A3(new_n570_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1336gat));
  OAI21_X1  g493(.A(G92gat), .B1(new_n692_), .B2(new_n297_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n297_), .A2(G92gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n688_), .B2(new_n696_), .ZN(G1337gat));
  OAI21_X1  g496(.A(G99gat), .B1(new_n692_), .B2(new_n383_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n609_), .A2(new_n467_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n698_), .B(new_n699_), .C1(new_n688_), .C2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT113), .Z(new_n703_));
  XNOR2_X1  g502(.A(new_n701_), .B(new_n703_), .ZN(G1338gat));
  NAND3_X1  g503(.A1(new_n625_), .A2(new_n342_), .A3(new_n691_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n468_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n707_), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n687_), .A2(new_n468_), .A3(new_n342_), .A4(new_n667_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n708_), .A2(new_n713_), .A3(new_n709_), .A4(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  INV_X1    g514(.A(KEYINPUT122), .ZN(new_n716_));
  INV_X1    g515(.A(G113gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n297_), .A2(new_n343_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n718_), .A2(new_n383_), .A3(new_n570_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n561_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n551_), .A2(new_n554_), .A3(new_n544_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT116), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n551_), .A2(new_n554_), .A3(KEYINPUT116), .A4(new_n544_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n539_), .A3(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n555_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(KEYINPUT55), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n728_), .B1(new_n555_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n720_), .B1(new_n725_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT56), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT117), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n556_), .A2(new_n561_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n734_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n720_), .B(new_n738_), .C1(new_n725_), .C2(new_n731_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n455_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT118), .B1(new_n737_), .B2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n739_), .A2(new_n455_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n732_), .A2(new_n734_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT118), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n443_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT119), .B(new_n451_), .C1(new_n446_), .C2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT119), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n438_), .B2(new_n445_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n453_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n438_), .A2(new_n441_), .A3(new_n746_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n454_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT120), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(KEYINPUT120), .A3(new_n454_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n563_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n741_), .A2(new_n745_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT57), .A3(new_n513_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT121), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT121), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(KEYINPUT57), .A4(new_n513_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n513_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n732_), .A2(KEYINPUT56), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n733_), .B(new_n720_), .C1(new_n725_), .C2(new_n731_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT58), .A3(new_n736_), .A4(new_n757_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n608_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n757_), .A2(new_n767_), .A3(new_n736_), .A4(new_n768_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT58), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n765_), .A2(new_n766_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n535_), .B1(new_n764_), .B2(new_n775_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n537_), .A2(new_n567_), .A3(new_n455_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT54), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n719_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n777_), .B(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n774_), .A2(new_n608_), .A3(new_n770_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n742_), .A2(new_n743_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n783_), .A2(KEYINPUT118), .B1(new_n563_), .B2(new_n757_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n574_), .B1(new_n784_), .B2(new_n745_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n785_), .B2(KEYINPUT57), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n781_), .B1(new_n787_), .B2(new_n536_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n719_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n779_), .A2(KEYINPUT59), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n717_), .B1(new_n791_), .B2(new_n455_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n779_), .A2(G113gat), .A3(new_n456_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n716_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n779_), .A2(KEYINPUT59), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n790_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n455_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G113gat), .ZN(new_n798_));
  INV_X1    g597(.A(new_n793_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(KEYINPUT122), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n794_), .A2(new_n800_), .ZN(G1340gat));
  INV_X1    g600(.A(new_n791_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G120gat), .B1(new_n802_), .B2(new_n576_), .ZN(new_n803_));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n576_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(KEYINPUT60), .B2(new_n804_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n779_), .B2(new_n806_), .ZN(G1341gat));
  INV_X1    g606(.A(new_n535_), .ZN(new_n808_));
  OAI21_X1  g607(.A(G127gat), .B1(new_n802_), .B2(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n598_), .A2(G127gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n779_), .B2(new_n810_), .ZN(G1342gat));
  OAI21_X1  g610(.A(G134gat), .B1(new_n802_), .B2(new_n514_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n513_), .A2(G134gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n779_), .B2(new_n813_), .ZN(G1343gat));
  NAND2_X1  g613(.A1(new_n764_), .A2(new_n775_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n808_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n781_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n297_), .A2(new_n383_), .A3(new_n342_), .A4(new_n370_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT123), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n456_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(new_n311_), .ZN(G1344gat));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n576_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(new_n312_), .ZN(G1345gat));
  NOR2_X1   g623(.A1(new_n820_), .A2(new_n598_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT61), .B(G155gat), .Z(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1346gat));
  INV_X1    g626(.A(new_n820_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G162gat), .B1(new_n828_), .B2(new_n574_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n608_), .A2(G162gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT124), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n828_), .B2(new_n831_), .ZN(G1347gat));
  NAND2_X1  g631(.A1(new_n585_), .A2(new_n384_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT125), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n342_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n536_), .B1(new_n764_), .B2(new_n775_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n455_), .B(new_n836_), .C1(new_n837_), .C2(new_n778_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G169gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n788_), .A2(new_n248_), .A3(new_n455_), .A4(new_n836_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT126), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n841_), .A2(new_n843_), .A3(KEYINPUT126), .A4(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1348gat));
  NAND2_X1  g647(.A1(new_n788_), .A2(new_n836_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G176gat), .B1(new_n850_), .B2(new_n567_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n342_), .B1(new_n816_), .B2(new_n781_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n835_), .A2(new_n576_), .A3(new_n249_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1349gat));
  NOR3_X1   g653(.A1(new_n849_), .A2(new_n240_), .A3(new_n808_), .ZN(new_n855_));
  INV_X1    g654(.A(G183gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(new_n536_), .A3(new_n834_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1350gat));
  OAI21_X1  g657(.A(G190gat), .B1(new_n849_), .B2(new_n514_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n574_), .A2(new_n241_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n849_), .B2(new_n860_), .ZN(G1351gat));
  NOR4_X1   g660(.A1(new_n297_), .A2(new_n609_), .A3(new_n343_), .A4(new_n370_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n817_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n456_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(new_n209_), .ZN(G1352gat));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n576_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(new_n207_), .ZN(G1353gat));
  NOR2_X1   g666(.A1(new_n863_), .A2(new_n808_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT63), .B(G211gat), .Z(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(new_n870_), .ZN(G1354gat));
  NOR3_X1   g670(.A1(new_n863_), .A2(new_n214_), .A3(new_n514_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n817_), .A2(new_n574_), .A3(new_n862_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT127), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G218gat), .B1(new_n873_), .B2(new_n874_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n872_), .B1(new_n875_), .B2(new_n876_), .ZN(G1355gat));
endmodule


