//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT10), .B(G99gat), .ZN(new_n206_));
  OAI221_X1 g005(.A(new_n204_), .B1(KEYINPUT9), .B2(new_n205_), .C1(G106gat), .C2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT64), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n202_), .A2(KEYINPUT8), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT65), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n212_), .B1(new_n210_), .B2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n216_), .A2(new_n209_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT8), .B1(new_n219_), .B2(new_n202_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n211_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT66), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n225_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G78gat), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT67), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n230_), .A2(KEYINPUT67), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n227_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n230_), .A2(KEYINPUT67), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n231_), .A3(new_n226_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n234_), .A2(KEYINPUT69), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT69), .B1(new_n234_), .B2(new_n236_), .ZN(new_n238_));
  OAI211_X1 g037(.A(KEYINPUT12), .B(new_n222_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n236_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n226_), .B1(new_n235_), .B2(new_n231_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n222_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT12), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n234_), .A2(new_n221_), .A3(new_n236_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G230gat), .A2(G233gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n234_), .A2(new_n236_), .A3(KEYINPUT68), .A4(new_n221_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n242_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n246_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT71), .ZN(new_n256_));
  XOR2_X1   g055(.A(G176gat), .B(G204gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  NAND3_X1  g059(.A1(new_n248_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT72), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n248_), .A2(new_n254_), .A3(new_n263_), .A4(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n248_), .A2(new_n254_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n265_), .A2(KEYINPUT13), .A3(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT13), .B1(new_n265_), .B2(new_n268_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G15gat), .B(G22gat), .Z(new_n272_));
  NAND2_X1  g071(.A1(G1gat), .A2(G8gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(KEYINPUT14), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT79), .ZN(new_n275_));
  XOR2_X1   g074(.A(G1gat), .B(G8gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G29gat), .B(G36gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT75), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G43gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G50gat), .ZN(new_n281_));
  INV_X1    g080(.A(G43gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n279_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G50gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT15), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n285_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT15), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n277_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G229gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n275_), .B(new_n276_), .Z(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(new_n288_), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n291_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G141gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G169gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(G197gat), .Z(new_n300_));
  NOR2_X1   g099(.A1(new_n286_), .A2(new_n277_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT81), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n295_), .B2(new_n301_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n297_), .B(new_n300_), .C1(new_n306_), .C2(new_n292_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n300_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n292_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(new_n296_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n271_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT104), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT86), .Z(new_n315_));
  XNOR2_X1  g114(.A(G15gat), .B(G43gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT82), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G169gat), .A3(G176gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT25), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G183gat), .ZN(new_n329_));
  INV_X1    g128(.A(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT26), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT26), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G190gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n327_), .A2(new_n329_), .A3(new_n331_), .A4(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n325_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n339_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n336_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G169gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT22), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT22), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G169gat), .ZN(new_n350_));
  INV_X1    g149(.A(G176gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT84), .B1(new_n337_), .B2(KEYINPUT23), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n355_), .A2(new_n344_), .A3(G183gat), .A4(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n341_), .A2(KEYINPUT23), .A3(new_n342_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n353_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n318_), .B1(new_n346_), .B2(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT83), .B1(G183gat), .B2(G190gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n344_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n338_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n367_), .A2(new_n325_), .A3(new_n335_), .A4(new_n334_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n360_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n368_), .B(KEYINPUT85), .C1(new_n369_), .C2(new_n353_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n371_), .A2(new_n372_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n317_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n317_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n315_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n315_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n376_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G134gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G127gat), .ZN(new_n384_));
  INV_X1    g183(.A(G127gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G134gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G120gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G113gat), .ZN(new_n389_));
  INV_X1    g188(.A(G113gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G120gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n384_), .A2(new_n386_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(KEYINPUT87), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n387_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT87), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n379_), .A2(new_n382_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n402_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT27), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT18), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G64gat), .ZN(new_n410_));
  INV_X1    g209(.A(G92gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n348_), .A2(new_n350_), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT97), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n351_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n322_), .A2(new_n324_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n367_), .A2(new_n361_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n359_), .A2(new_n335_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n332_), .A2(G190gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n330_), .A2(KEYINPUT26), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n327_), .A2(new_n329_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n331_), .A2(new_n333_), .A3(KEYINPUT94), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n320_), .A2(new_n321_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n429_), .A2(KEYINPUT95), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT95), .B1(new_n429_), .B2(new_n430_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n422_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT96), .B(new_n422_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n420_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G197gat), .B(G204gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(G211gat), .B(G218gat), .Z(new_n439_));
  INV_X1    g238(.A(KEYINPUT21), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n439_), .A2(new_n440_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n437_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G226gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT19), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n363_), .A2(new_n370_), .A3(new_n443_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT20), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT93), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n453_), .A3(KEYINPUT20), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n452_), .B(new_n454_), .C1(new_n443_), .C2(new_n437_), .ZN(new_n455_));
  AOI221_X4 g254(.A(new_n413_), .B1(new_n444_), .B2(new_n449_), .C1(new_n455_), .C2(new_n448_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n448_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n444_), .A2(new_n449_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n412_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n407_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT90), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT90), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT2), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n465_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G155gat), .ZN(new_n475_));
  INV_X1    g274(.A(G162gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G155gat), .A2(G162gat), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G141gat), .B(G148gat), .Z(new_n481_));
  INV_X1    g280(.A(KEYINPUT88), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n478_), .A2(new_n482_), .A3(KEYINPUT1), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n478_), .B2(KEYINPUT1), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT89), .B1(new_n478_), .B2(KEYINPUT1), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT1), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(G155gat), .A4(G162gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n489_), .A3(new_n477_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n481_), .B1(new_n485_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n480_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n443_), .B1(KEYINPUT29), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G78gat), .B(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n493_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT91), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n443_), .B2(KEYINPUT92), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n496_), .B(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n492_), .A2(KEYINPUT29), .ZN(new_n501_));
  XOR2_X1   g300(.A(G22gat), .B(G50gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT28), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n501_), .B(new_n503_), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n496_), .A2(new_n499_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n496_), .A2(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n412_), .B(KEYINPUT103), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n455_), .A2(new_n448_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n448_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n443_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n419_), .A2(new_n433_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(KEYINPUT100), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(KEYINPUT100), .B2(new_n515_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n445_), .A2(new_n446_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n513_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n511_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n457_), .A2(new_n458_), .A3(new_n412_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(KEYINPUT27), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n460_), .A2(new_n510_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n393_), .A2(new_n394_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n480_), .A2(new_n491_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n488_), .A2(G155gat), .A3(G162gat), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n526_), .A2(KEYINPUT89), .B1(new_n475_), .B2(new_n476_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n527_), .B(new_n489_), .C1(new_n484_), .C2(new_n483_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n528_), .A2(new_n481_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n395_), .A2(new_n398_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n525_), .B(KEYINPUT4), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT98), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n492_), .A2(new_n399_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT98), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT4), .A4(new_n525_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n529_), .A2(new_n530_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G225gat), .A2(G233gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT99), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G1gat), .B(G29gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT0), .ZN(new_n544_));
  INV_X1    g343(.A(G57gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(G85gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n533_), .A2(new_n525_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n541_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n542_), .A2(KEYINPUT101), .A3(new_n548_), .A4(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n548_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n531_), .A2(KEYINPUT98), .B1(new_n536_), .B2(new_n537_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n550_), .B1(new_n557_), .B2(new_n535_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n551_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n556_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT102), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n554_), .A2(KEYINPUT102), .A3(new_n555_), .A4(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n523_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n429_), .A2(new_n430_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n429_), .A2(KEYINPUT95), .A3(new_n430_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT96), .B1(new_n571_), .B2(new_n422_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n436_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n419_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n574_), .A2(new_n514_), .B1(KEYINPUT93), .B2(new_n451_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n513_), .B1(new_n575_), .B2(new_n454_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n458_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n413_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n539_), .A2(new_n541_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n560_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n560_), .A2(new_n582_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n578_), .A2(new_n583_), .A3(new_n584_), .A4(new_n521_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n457_), .A2(new_n458_), .A3(new_n586_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n561_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n510_), .B1(new_n585_), .B2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n313_), .B(new_n406_), .C1(new_n566_), .C2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n510_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n460_), .A3(new_n522_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n594_), .A2(new_n406_), .A3(new_n565_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n406_), .B1(new_n566_), .B2(new_n591_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n596_), .B2(KEYINPUT104), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n312_), .B1(new_n592_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT73), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT34), .ZN(new_n603_));
  OAI22_X1  g402(.A1(new_n222_), .A2(new_n288_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n287_), .A2(new_n290_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n605_), .B2(new_n222_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n600_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n221_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n600_), .B(new_n603_), .C1(new_n609_), .C2(new_n604_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n610_), .A3(KEYINPUT78), .ZN(new_n611_));
  XOR2_X1   g410(.A(G134gat), .B(G162gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  NAND2_X1  g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n608_), .A2(new_n610_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n611_), .A2(new_n620_), .A3(new_n616_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT17), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT16), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n326_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n277_), .B(KEYINPUT80), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n237_), .A2(new_n238_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n629_), .B(new_n633_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n637_), .B2(new_n636_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n633_), .B(new_n629_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n240_), .A2(new_n241_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n641_), .B2(new_n636_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n628_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n598_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT105), .ZN(new_n647_));
  INV_X1    g446(.A(new_n565_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(G1gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(KEYINPUT38), .A3(new_n649_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n622_), .A2(new_n654_), .A3(new_n624_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n644_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n598_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G1gat), .B1(new_n660_), .B2(new_n648_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n652_), .A2(new_n653_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n652_), .A2(KEYINPUT107), .A3(new_n653_), .A4(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1324gat));
  INV_X1    g465(.A(G8gat), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n460_), .A2(new_n522_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n647_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n660_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n669_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(G8gat), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n672_), .B2(G8gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n670_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n647_), .A2(new_n679_), .A3(new_n405_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n671_), .A2(new_n405_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n681_), .B2(G15gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT109), .ZN(G1326gat));
  OAI21_X1  g484(.A(G22gat), .B1(new_n660_), .B2(new_n593_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT42), .ZN(new_n687_));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n647_), .A2(new_n688_), .A3(new_n510_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1327gat));
  INV_X1    g489(.A(new_n644_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n691_), .B(new_n657_), .C1(new_n597_), .C2(new_n592_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n312_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n565_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n312_), .A2(new_n691_), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT43), .B(new_n627_), .C1(new_n597_), .C2(new_n592_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n460_), .A2(new_n510_), .A3(new_n522_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n591_), .B1(new_n700_), .B2(new_n648_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT104), .B1(new_n701_), .B2(new_n405_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n595_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n592_), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n699_), .B1(new_n704_), .B2(new_n628_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n697_), .B1(new_n698_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n697_), .C1(new_n698_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n565_), .A2(G29gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n696_), .B1(new_n711_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n668_), .A2(G36gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n692_), .A2(new_n693_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT45), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n692_), .A2(new_n720_), .A3(new_n693_), .A4(new_n717_), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n719_), .A2(new_n721_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n708_), .A2(new_n669_), .A3(new_n709_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(KEYINPUT110), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n708_), .A2(new_n727_), .A3(new_n669_), .A4(new_n709_), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n716_), .B(new_n723_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n716_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n725_), .A2(KEYINPUT110), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(G36gat), .A3(new_n728_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n732_), .B2(new_n722_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n729_), .A2(new_n733_), .ZN(G1329gat));
  NOR3_X1   g533(.A1(new_n694_), .A2(G43gat), .A3(new_n406_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n708_), .A2(new_n405_), .A3(new_n709_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G43gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g537(.A(G50gat), .B1(new_n710_), .B2(new_n593_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n510_), .A2(new_n284_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT112), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n694_), .B2(new_n741_), .ZN(G1331gat));
  NOR2_X1   g541(.A1(new_n271_), .A2(new_n311_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n704_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n645_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n545_), .A3(new_n565_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(KEYINPUT113), .A3(new_n659_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n659_), .A2(new_n704_), .A3(new_n743_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n565_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n747_), .B1(new_n753_), .B2(new_n545_), .ZN(G1332gat));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n746_), .A2(new_n755_), .A3(new_n669_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n752_), .A2(new_n669_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G64gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT48), .B(new_n755_), .C1(new_n752_), .C2(new_n669_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1333gat));
  OR3_X1    g560(.A1(new_n745_), .A2(G71gat), .A3(new_n406_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n748_), .A2(new_n405_), .A3(new_n751_), .ZN(new_n763_));
  XOR2_X1   g562(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(G71gat), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G71gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT115), .ZN(G1334gat));
  INV_X1    g567(.A(G78gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n746_), .A2(new_n769_), .A3(new_n510_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n752_), .A2(new_n510_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G78gat), .ZN(new_n773_));
  AOI211_X1 g572(.A(KEYINPUT50), .B(new_n769_), .C1(new_n752_), .C2(new_n510_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1335gat));
  NAND2_X1  g574(.A1(new_n743_), .A2(new_n644_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n698_), .A2(new_n705_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n778_), .B2(new_n777_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780_), .B2(new_n648_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n692_), .A2(new_n743_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n547_), .A3(new_n565_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n780_), .B2(new_n668_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n411_), .A3(new_n669_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n780_), .B2(new_n406_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n406_), .A2(new_n206_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n782_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT51), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n788_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n743_), .A2(new_n510_), .A3(new_n644_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n777_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  INV_X1    g599(.A(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT117), .B1(new_n797_), .B2(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n800_), .A2(KEYINPUT52), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n782_), .A2(new_n801_), .A3(new_n510_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n802_), .B2(KEYINPUT52), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(KEYINPUT52), .A3(new_n802_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n802_), .A2(KEYINPUT52), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .A4(new_n804_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(G1339gat));
  NAND2_X1  g610(.A1(new_n622_), .A2(new_n624_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT37), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n311_), .B1(new_n814_), .B2(KEYINPUT54), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n816_));
  AND4_X1   g615(.A1(new_n691_), .A2(new_n813_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n817_), .B(new_n271_), .C1(new_n814_), .C2(KEYINPUT54), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n627_), .A2(new_n691_), .A3(new_n815_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n271_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n265_), .A2(new_n311_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n239_), .A2(new_n250_), .A3(new_n244_), .A4(new_n251_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n253_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n239_), .A2(KEYINPUT55), .A3(new_n244_), .A4(new_n247_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n248_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n267_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n267_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n824_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n303_), .A2(new_n305_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n292_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n291_), .A2(new_n838_), .A3(new_n295_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n291_), .B2(new_n295_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n293_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n837_), .B(new_n308_), .C1(new_n839_), .C2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n307_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n657_), .B(KEYINPUT57), .C1(new_n835_), .C2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n267_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n267_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n265_), .A2(new_n268_), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n850_), .A2(new_n824_), .B1(new_n851_), .B2(new_n843_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n657_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n833_), .A2(new_n834_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n824_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n844_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n854_), .B1(new_n857_), .B2(new_n658_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  INV_X1    g658(.A(new_n843_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n265_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n859_), .B1(new_n850_), .B2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n855_), .A2(KEYINPUT58), .A3(new_n265_), .A4(new_n860_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n628_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n847_), .A2(new_n853_), .A3(new_n858_), .A4(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n823_), .B1(new_n865_), .B2(new_n644_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n594_), .A2(new_n648_), .A3(new_n406_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n390_), .A3(new_n311_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n311_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n865_), .A2(new_n644_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n823_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n875_), .B2(new_n867_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n866_), .A2(new_n868_), .A3(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT122), .B1(new_n876_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT59), .B1(new_n866_), .B2(new_n868_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n875_), .A2(new_n867_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n881_), .B(new_n882_), .C1(new_n883_), .C2(new_n878_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n871_), .B1(new_n880_), .B2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n870_), .B1(new_n885_), .B2(new_n390_), .ZN(G1340gat));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n271_), .B2(G120gat), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n869_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n887_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n889_), .A2(new_n876_), .A3(new_n271_), .A4(new_n879_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n388_), .ZN(G1341gat));
  NAND3_X1  g691(.A1(new_n869_), .A2(new_n385_), .A3(new_n691_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n644_), .B1(new_n880_), .B2(new_n884_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n385_), .ZN(G1342gat));
  NAND3_X1  g694(.A1(new_n869_), .A2(new_n383_), .A3(new_n658_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n627_), .B1(new_n880_), .B2(new_n884_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n383_), .ZN(G1343gat));
  NOR3_X1   g697(.A1(new_n648_), .A2(new_n523_), .A3(new_n405_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n875_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n871_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n471_), .ZN(G1344gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n271_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n472_), .ZN(G1345gat));
  NOR2_X1   g703(.A1(new_n900_), .A2(new_n644_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT61), .B(G155gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n900_), .B2(new_n627_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n658_), .A2(new_n476_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n900_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT123), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n908_), .B(new_n912_), .C1(new_n900_), .C2(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1347gat));
  NAND4_X1  g713(.A1(new_n669_), .A2(new_n405_), .A3(new_n593_), .A4(new_n648_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n866_), .A2(new_n871_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  OAI21_X1  g716(.A(G169gat), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n917_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n919_), .A2(KEYINPUT62), .A3(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  INV_X1    g721(.A(new_n920_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n918_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n916_), .A2(new_n415_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n921_), .A2(new_n924_), .A3(new_n925_), .ZN(G1348gat));
  XNOR2_X1  g725(.A(KEYINPUT125), .B(G176gat), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n351_), .A2(KEYINPUT125), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n866_), .A2(new_n915_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n821_), .ZN(new_n930_));
  MUX2_X1   g729(.A(new_n927_), .B(new_n928_), .S(new_n930_), .Z(G1349gat));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  AOI21_X1  g731(.A(G183gat), .B1(new_n929_), .B2(new_n691_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n427_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n929_), .A2(new_n935_), .A3(new_n691_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n932_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n936_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n938_), .A2(KEYINPUT126), .A3(new_n933_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1350gat));
  AOI21_X1  g739(.A(new_n330_), .B1(new_n929_), .B2(new_n628_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n929_), .A2(new_n426_), .A3(new_n428_), .A4(new_n658_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1351gat));
  NAND3_X1  g743(.A1(new_n669_), .A2(new_n406_), .A3(new_n510_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n866_), .A2(new_n565_), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n311_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n821_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g749(.A1(new_n946_), .A2(new_n691_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AND2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  INV_X1    g754(.A(G218gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n946_), .A2(new_n956_), .A3(new_n658_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n946_), .A2(new_n628_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n956_), .ZN(G1355gat));
endmodule


