//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT81), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(KEYINPUT23), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(KEYINPUT81), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT78), .B(G183gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n212_), .B(KEYINPUT80), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(new_n209_), .B2(KEYINPUT25), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT26), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n223_), .A2(KEYINPUT79), .A3(KEYINPUT26), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT79), .B1(new_n223_), .B2(KEYINPUT26), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n207_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n211_), .B1(new_n220_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT82), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n211_), .B(KEYINPUT82), .C1(new_n220_), .C2(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G43gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT30), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G15gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n235_), .A2(new_n240_), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT84), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT84), .B1(new_n241_), .B2(new_n242_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  INV_X1    g044(.A(G113gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G120gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n244_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n244_), .A2(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G64gat), .B(G92gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G8gat), .B(G36gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  INV_X1    g060(.A(KEYINPUT96), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263_));
  INV_X1    g062(.A(G197gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(G204gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(G204gat), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(KEYINPUT90), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n267_), .A2(KEYINPUT91), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n269_), .B(new_n268_), .C1(new_n266_), .C2(new_n265_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT91), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274_));
  INV_X1    g073(.A(new_n266_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n264_), .A2(G204gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(KEYINPUT21), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n270_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n267_), .A2(new_n269_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n268_), .B1(new_n274_), .B2(KEYINPUT92), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n280_), .B(new_n281_), .C1(KEYINPUT92), .C2(new_n274_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n231_), .A2(new_n283_), .A3(new_n232_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n282_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT95), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n215_), .A2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n287_), .B(new_n289_), .C1(new_n288_), .C2(new_n203_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n223_), .A2(KEYINPUT26), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n224_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT25), .B(G183gat), .Z(new_n293_));
  OAI221_X1 g092(.A(new_n206_), .B1(new_n292_), .B2(new_n293_), .C1(KEYINPUT81), .C2(new_n207_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n294_), .B2(new_n220_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n285_), .B1(new_n286_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n284_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G226gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT19), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT94), .Z(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n262_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  AOI211_X1 g101(.A(KEYINPUT96), .B(new_n300_), .C1(new_n284_), .C2(new_n296_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n285_), .B1(new_n233_), .B2(new_n286_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n299_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n286_), .A2(new_n295_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n261_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n297_), .A2(new_n301_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT96), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n297_), .A2(new_n262_), .A3(new_n301_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n312_), .A2(new_n261_), .A3(new_n309_), .A4(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n256_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n261_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n306_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n297_), .A2(new_n301_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(KEYINPUT27), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT102), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  INV_X1    g123(.A(G155gat), .ZN(new_n325_));
  INV_X1    g124(.A(G162gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n327_), .B(new_n328_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT88), .ZN(new_n330_));
  OR2_X1    g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n331_), .A2(KEYINPUT3), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(KEYINPUT3), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n332_), .A2(new_n335_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(KEYINPUT88), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n330_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n331_), .B(KEYINPUT85), .ZN(new_n341_));
  AND3_X1   g140(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n327_), .B(new_n328_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n333_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n341_), .A2(KEYINPUT87), .A3(new_n333_), .A4(new_n344_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n340_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n349_), .A2(KEYINPUT29), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT28), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(KEYINPUT28), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G50gat), .ZN(new_n354_));
  INV_X1    g153(.A(G50gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n355_), .A3(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n349_), .A2(KEYINPUT29), .ZN(new_n358_));
  AND2_X1   g157(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(G233gat), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n361_), .A3(new_n286_), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n363_));
  AOI21_X1  g162(.A(new_n283_), .B1(new_n349_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n364_), .B2(new_n361_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366_));
  INV_X1    g165(.A(G22gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n362_), .B(new_n370_), .C1(new_n364_), .C2(new_n361_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n357_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n354_), .A2(new_n369_), .A3(new_n356_), .A4(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n283_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n376_), .A2(new_n285_), .A3(new_n307_), .ZN(new_n377_));
  OAI22_X1  g176(.A1(new_n377_), .A2(new_n306_), .B1(new_n301_), .B2(new_n297_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n256_), .B1(new_n378_), .B2(new_n317_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT102), .A3(new_n314_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n316_), .A2(new_n323_), .A3(new_n375_), .A4(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n347_), .A2(new_n348_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT98), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n249_), .A4(new_n340_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n247_), .B(G120gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n349_), .B2(KEYINPUT98), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(new_n386_), .A3(KEYINPUT4), .ZN(new_n390_));
  INV_X1    g189(.A(new_n388_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(KEYINPUT99), .A2(KEYINPUT4), .ZN(new_n392_));
  AND2_X1   g191(.A1(KEYINPUT99), .A2(KEYINPUT4), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n349_), .B(new_n385_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT100), .B(KEYINPUT0), .Z(new_n397_));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G57gat), .B(G85gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n396_), .B(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n381_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n378_), .A2(KEYINPUT32), .A3(new_n261_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n261_), .A2(KEYINPUT32), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n312_), .A2(new_n309_), .A3(new_n313_), .A4(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n407_), .A2(KEYINPUT101), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(KEYINPUT101), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n403_), .B(new_n405_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n389_), .A2(new_n395_), .A3(new_n402_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT33), .ZN(new_n412_));
  INV_X1    g211(.A(new_n310_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n387_), .A2(new_n391_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n390_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n401_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n412_), .A2(new_n413_), .A3(new_n314_), .A4(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n375_), .B1(new_n410_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n255_), .B1(new_n404_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n374_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n354_), .A2(new_n356_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n316_), .A2(new_n422_), .A3(new_n323_), .A4(new_n380_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT103), .ZN(new_n424_));
  AND4_X1   g223(.A1(KEYINPUT102), .A2(new_n314_), .A3(KEYINPUT27), .A4(new_n320_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT102), .B1(new_n379_), .B2(new_n314_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT103), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n422_), .A4(new_n316_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n403_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n255_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n424_), .A2(new_n429_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n419_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT71), .ZN(new_n434_));
  INV_X1    g233(.A(G71gat), .ZN(new_n435_));
  INV_X1    g234(.A(G78gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n436_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G57gat), .B(G64gat), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n438_), .B(new_n439_), .C1(new_n440_), .C2(KEYINPUT11), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT70), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n440_), .B2(KEYINPUT11), .ZN(new_n443_));
  AND2_X1   g242(.A1(G57gat), .A2(G64gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G57gat), .A2(G64gat), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n442_), .B(KEYINPUT11), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n441_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n444_), .A2(new_n445_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT11), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n437_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT11), .B1(new_n444_), .B2(new_n445_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT70), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n439_), .A2(new_n451_), .B1(new_n453_), .B2(new_n446_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n434_), .B1(new_n448_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n441_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n451_), .A2(new_n453_), .A3(new_n446_), .A4(new_n439_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT71), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT10), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT10), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G99gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT66), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G99gat), .A3(G106gat), .ZN(new_n474_));
  AND2_X1   g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT9), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n472_), .A2(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(KEYINPUT67), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT9), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G85gat), .A2(G92gat), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n479_), .A2(new_n480_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n470_), .A2(new_n477_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n470_), .A2(new_n477_), .A3(new_n484_), .A4(KEYINPUT68), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n475_), .A2(new_n478_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n472_), .A2(new_n474_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n490_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT8), .B1(new_n490_), .B2(KEYINPUT69), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n497_), .B(new_n490_), .C1(new_n491_), .C2(new_n495_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT12), .B1(new_n459_), .B2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n455_), .A2(new_n458_), .A3(new_n501_), .A4(new_n489_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G230gat), .A2(G233gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT64), .Z(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT65), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n456_), .A2(new_n457_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(KEYINPUT12), .A3(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n455_), .A2(new_n458_), .B1(new_n501_), .B2(new_n489_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n509_), .B1(new_n505_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G120gat), .B(G148gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G176gat), .ZN(new_n518_));
  INV_X1    g317(.A(G204gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n515_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G29gat), .B(G36gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G43gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(new_n355_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n532_), .B(new_n234_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(G50gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n531_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(G50gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(new_n355_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(KEYINPUT15), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542_));
  INV_X1    g341(.A(G1gat), .ZN(new_n543_));
  INV_X1    g342(.A(G8gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT14), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G1gat), .B(G8gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n541_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n534_), .A2(new_n536_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n548_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT76), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n538_), .A2(new_n539_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n551_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n549_), .A2(new_n556_), .A3(KEYINPUT76), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563_));
  INV_X1    g362(.A(G169gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n264_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n554_), .A2(new_n561_), .A3(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n567_), .A2(KEYINPUT77), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT77), .B1(new_n567_), .B2(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n530_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n541_), .A2(new_n502_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n552_), .A2(new_n501_), .A3(new_n489_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT35), .Z(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(new_n576_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT73), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n575_), .A2(KEYINPUT73), .A3(new_n576_), .A4(new_n579_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G134gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n326_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n575_), .A2(new_n576_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(KEYINPUT35), .A3(new_n578_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n584_), .A2(new_n585_), .A3(new_n588_), .A4(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n585_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n588_), .A2(new_n585_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n591_), .A2(new_n592_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n548_), .B(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(new_n511_), .Z(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n602_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n459_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n612_), .B2(new_n601_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n609_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n613_), .B(new_n614_), .C1(new_n612_), .C2(new_n601_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT37), .A4(new_n596_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n599_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n433_), .A2(new_n574_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT104), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n543_), .A3(new_n403_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n433_), .A2(new_n574_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n591_), .A2(new_n596_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT105), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n624_), .A2(new_n625_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n430_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n621_), .A2(new_n622_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n623_), .A2(new_n631_), .A3(new_n632_), .ZN(G1324gat));
  NAND2_X1  g432(.A1(new_n427_), .A2(new_n316_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n620_), .A2(new_n544_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n629_), .A2(new_n634_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(G8gat), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT39), .B(new_n544_), .C1(new_n629_), .C2(new_n634_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n630_), .B2(new_n255_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT41), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n619_), .A2(G15gat), .A3(new_n255_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  AOI21_X1  g444(.A(new_n367_), .B1(new_n629_), .B2(new_n375_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT42), .Z(new_n647_));
  NAND2_X1  g446(.A1(new_n375_), .A2(new_n367_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n619_), .B2(new_n648_), .ZN(G1327gat));
  NOR3_X1   g448(.A1(new_n624_), .A2(new_n616_), .A3(new_n626_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n403_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n599_), .A2(new_n617_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n433_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT107), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n433_), .A2(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n433_), .A2(new_n659_), .A3(new_n652_), .A4(new_n654_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n574_), .A2(new_n625_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT106), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n663_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n664_), .A2(G29gat), .A3(new_n403_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n663_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n651_), .B1(new_n665_), .B2(new_n668_), .ZN(G1328gat));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n634_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n671_), .B1(new_n673_), .B2(new_n664_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n650_), .A2(new_n671_), .A3(new_n634_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n670_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n664_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT44), .B1(new_n661_), .B2(new_n663_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n672_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT46), .B(new_n676_), .C1(new_n681_), .C2(new_n671_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n678_), .A2(new_n682_), .ZN(G1329gat));
  NAND4_X1  g482(.A1(new_n668_), .A2(G43gat), .A3(new_n431_), .A4(new_n664_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n650_), .A2(new_n431_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n234_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n684_), .A2(new_n688_), .A3(new_n686_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1330gat));
  AOI21_X1  g491(.A(G50gat), .B1(new_n650_), .B2(new_n375_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n680_), .A2(new_n355_), .A3(new_n422_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n664_), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n529_), .A2(new_n572_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n433_), .A2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(new_n618_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n403_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n433_), .A2(new_n616_), .A3(new_n627_), .A4(new_n696_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n403_), .A2(G57gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(G1332gat));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n700_), .B2(new_n634_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT48), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n634_), .A2(new_n703_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT109), .Z(new_n707_));
  NAND2_X1  g506(.A1(new_n698_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1333gat));
  AOI21_X1  g508(.A(new_n435_), .B1(new_n700_), .B2(new_n431_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT49), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n698_), .A2(new_n435_), .A3(new_n431_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1334gat));
  NAND3_X1  g512(.A1(new_n698_), .A2(new_n436_), .A3(new_n375_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n700_), .A2(new_n375_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G78gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n717_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1335gat));
  AND4_X1   g521(.A1(new_n625_), .A2(new_n697_), .A3(new_n591_), .A4(new_n596_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n403_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n529_), .A2(new_n572_), .A3(new_n616_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n661_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n403_), .A2(G85gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1336gat));
  AOI21_X1  g528(.A(G92gat), .B1(new_n723_), .B2(new_n634_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n634_), .A2(G92gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT112), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n727_), .B2(new_n732_), .ZN(G1337gat));
  OAI21_X1  g532(.A(G99gat), .B1(new_n726_), .B2(new_n255_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n723_), .A2(new_n464_), .A3(new_n431_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT114), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n734_), .A2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT51), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT114), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n734_), .A2(new_n741_), .A3(new_n735_), .A4(new_n736_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(new_n740_), .A3(new_n742_), .ZN(G1338gat));
  NAND3_X1  g542(.A1(new_n723_), .A2(new_n469_), .A3(new_n375_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n661_), .A2(new_n375_), .A3(new_n725_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G106gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n744_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1339gat));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n618_), .A2(new_n754_), .A3(new_n573_), .A4(new_n529_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n599_), .A2(new_n573_), .A3(new_n616_), .A4(new_n617_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT115), .B1(new_n756_), .B2(new_n530_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n757_), .A3(KEYINPUT54), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n512_), .B(new_n504_), .C1(new_n514_), .C2(KEYINPUT12), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n509_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OR2_X1    g565(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n506_), .A2(new_n510_), .A3(new_n512_), .A4(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n763_), .B2(new_n509_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n763_), .A2(KEYINPUT117), .A3(new_n509_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n766_), .A2(new_n768_), .A3(new_n770_), .A4(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n520_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT56), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n550_), .A2(new_n559_), .A3(new_n553_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n558_), .A2(new_n551_), .A3(new_n560_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n566_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n569_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n772_), .A2(new_n779_), .A3(new_n520_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n774_), .A2(new_n522_), .A3(new_n778_), .A4(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT118), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT58), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT118), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n654_), .A3(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n774_), .A2(new_n572_), .A3(new_n522_), .A4(new_n780_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n778_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT57), .A3(new_n626_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n626_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n786_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n625_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n762_), .A2(new_n795_), .ZN(new_n796_));
  AND4_X1   g595(.A1(new_n403_), .A2(new_n424_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n572_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n755_), .A2(KEYINPUT54), .A3(new_n757_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT54), .B1(new_n755_), .B2(new_n757_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n781_), .A2(KEYINPUT118), .A3(new_n784_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n784_), .B1(new_n781_), .B2(KEYINPUT118), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n653_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n789_), .B2(new_n626_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n786_), .A2(KEYINPUT119), .A3(new_n793_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n790_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n803_), .B1(new_n811_), .B2(new_n625_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n797_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(KEYINPUT59), .B2(new_n798_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n573_), .A2(new_n246_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n800_), .B1(new_n816_), .B2(new_n817_), .ZN(G1340gat));
  OAI21_X1  g617(.A(new_n248_), .B1(new_n529_), .B2(KEYINPUT60), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n799_), .B(new_n819_), .C1(KEYINPUT60), .C2(new_n248_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n816_), .A2(new_n530_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n248_), .ZN(G1341gat));
  AOI21_X1  g621(.A(G127gat), .B1(new_n799_), .B2(new_n616_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n616_), .A2(G127gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n816_), .B2(new_n824_), .ZN(G1342gat));
  INV_X1    g624(.A(G134gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n798_), .B2(new_n627_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n653_), .A2(new_n826_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n828_), .B(new_n829_), .C1(new_n816_), .C2(new_n830_), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n796_), .A2(new_n255_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(new_n430_), .A3(new_n381_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n572_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n530_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n616_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT61), .B(G155gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1346gat));
  AOI21_X1  g639(.A(G162gat), .B1(new_n833_), .B2(new_n628_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n653_), .A2(new_n326_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n833_), .B2(new_n842_), .ZN(G1347gat));
  NAND2_X1  g642(.A1(new_n810_), .A2(new_n790_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT119), .B1(new_n786_), .B2(new_n793_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n625_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n375_), .B1(new_n846_), .B2(new_n762_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n672_), .A2(new_n403_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n255_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT22), .B(G169gat), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n847_), .A2(new_n572_), .A3(new_n850_), .A4(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n572_), .A3(new_n431_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT121), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT122), .B1(new_n847_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n812_), .A2(new_n858_), .A3(new_n375_), .A4(new_n855_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n853_), .B1(new_n860_), .B2(G169gat), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n857_), .A2(new_n859_), .A3(KEYINPUT62), .A4(new_n564_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n852_), .B1(new_n861_), .B2(new_n862_), .ZN(G1348gat));
  AND2_X1   g662(.A1(new_n847_), .A2(new_n850_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G176gat), .B1(new_n864_), .B2(new_n530_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n796_), .A2(KEYINPUT123), .A3(new_n422_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n760_), .A2(new_n761_), .B1(new_n794_), .B2(new_n625_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n375_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n866_), .A2(new_n869_), .A3(new_n850_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n530_), .A2(G176gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n865_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  AND3_X1   g671(.A1(new_n864_), .A2(new_n293_), .A3(new_n616_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n866_), .A2(new_n869_), .A3(new_n616_), .A4(new_n850_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT124), .ZN(new_n875_));
  INV_X1    g674(.A(new_n209_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n875_), .B2(new_n876_), .ZN(G1350gat));
  NAND4_X1  g676(.A1(new_n864_), .A2(new_n291_), .A3(new_n224_), .A4(new_n628_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n864_), .A2(new_n654_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n223_), .ZN(G1351gat));
  NAND4_X1  g679(.A1(new_n796_), .A2(new_n375_), .A3(new_n255_), .A4(new_n848_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n573_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(new_n264_), .ZN(G1352gat));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n529_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n519_), .ZN(G1353gat));
  INV_X1    g684(.A(new_n881_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n887_));
  INV_X1    g686(.A(G211gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n886_), .A2(new_n616_), .A3(new_n889_), .A4(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n887_), .B(new_n888_), .C1(new_n881_), .C2(new_n625_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1354gat));
  NAND3_X1  g694(.A1(new_n886_), .A2(KEYINPUT127), .A3(new_n628_), .ZN(new_n896_));
  INV_X1    g695(.A(G218gat), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n881_), .B2(new_n627_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n897_), .A3(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n886_), .A2(G218gat), .A3(new_n654_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1355gat));
endmodule


