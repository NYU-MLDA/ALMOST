//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G29gat), .B(G36gat), .Z(new_n208_));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209_));
  XOR2_X1   g008(.A(new_n208_), .B(new_n209_), .Z(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT15), .Z(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(new_n223_), .B2(KEYINPUT65), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n219_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(new_n217_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n223_), .B1(new_n231_), .B2(new_n216_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n227_), .ZN(new_n233_));
  OR2_X1    g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n221_), .A2(KEYINPUT9), .A3(new_n222_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n222_), .A2(KEYINPUT9), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n216_), .A4(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n229_), .A2(new_n233_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n211_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n232_), .B2(new_n227_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n227_), .A2(new_n220_), .A3(new_n224_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n229_), .A2(new_n233_), .A3(new_n246_), .A4(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n242_), .B1(new_n248_), .B2(new_n210_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(KEYINPUT69), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT35), .ZN(new_n252_));
  XOR2_X1   g051(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT35), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n249_), .A2(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n250_), .A2(new_n254_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n207_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n205_), .B(KEYINPUT36), .Z(new_n261_));
  AND4_X1   g060(.A1(new_n259_), .A2(new_n257_), .A3(new_n255_), .A4(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n202_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT71), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268_));
  INV_X1    g067(.A(G43gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(G15gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n270_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT23), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT81), .B(G190gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n276_), .B1(G183gat), .B2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G169gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n277_), .B2(KEYINPUT26), .ZN(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT25), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n284_), .A2(KEYINPUT25), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n283_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT24), .A3(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n276_), .B(new_n295_), .C1(KEYINPUT24), .C2(new_n293_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n281_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT82), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT84), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n274_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n301_), .B2(new_n300_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n274_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT85), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G113gat), .B(G120gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n307_), .A2(KEYINPUT85), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(KEYINPUT85), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n309_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT31), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n305_), .A2(new_n306_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n305_), .A2(new_n306_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n316_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n305_), .A2(new_n306_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n317_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n324_), .B2(KEYINPUT1), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n325_), .B2(KEYINPUT87), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(KEYINPUT87), .B2(new_n325_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  OR2_X1    g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n324_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n328_), .B(KEYINPUT2), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(new_n329_), .B2(KEYINPUT88), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n329_), .A2(KEYINPUT88), .A3(KEYINPUT3), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n322_), .B(new_n331_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT28), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(KEYINPUT28), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G22gat), .B(G50gat), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G211gat), .B(G218gat), .Z(new_n347_));
  INV_X1    g146(.A(KEYINPUT21), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G197gat), .B(G204gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n349_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n347_), .A3(KEYINPUT21), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n346_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G228gat), .A3(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT92), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT93), .Z(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n354_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G228gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT89), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n356_), .A2(new_n357_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n358_), .A2(new_n360_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n358_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n360_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT95), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n344_), .B(new_n369_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT95), .B1(new_n370_), .B2(new_n371_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI211_X1 g175(.A(KEYINPUT94), .B(new_n344_), .C1(new_n372_), .C2(new_n369_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT94), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n369_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n344_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OR3_X1    g180(.A1(new_n376_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(KEYINPUT97), .Z(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(G169gat), .B2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT99), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n292_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n389_), .B2(new_n388_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(new_n285_), .A3(new_n289_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n292_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n393_), .A2(new_n276_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n276_), .B1(G183gat), .B2(G190gat), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT100), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(KEYINPUT100), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n280_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n354_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT101), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT101), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n404_), .A3(new_n354_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n298_), .B2(new_n362_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n386_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n298_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n407_), .B1(new_n411_), .B2(new_n363_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n401_), .A2(new_n354_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(new_n385_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT18), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n410_), .A2(new_n415_), .A3(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n406_), .A2(new_n408_), .A3(new_n386_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n385_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n354_), .B1(new_n401_), .B2(KEYINPUT105), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(KEYINPUT105), .B2(new_n401_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n412_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n421_), .B1(new_n427_), .B2(new_n420_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G85gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n337_), .A2(new_n315_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n436_), .B2(KEYINPUT4), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n311_), .A2(new_n314_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n330_), .A3(new_n336_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(KEYINPUT4), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT102), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT102), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n436_), .A2(new_n442_), .A3(KEYINPUT4), .A4(new_n439_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT103), .B(new_n437_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n436_), .A2(new_n439_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(new_n435_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n437_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT103), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n433_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n450_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n432_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n428_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n410_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n441_), .A2(new_n443_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n456_), .B(new_n434_), .C1(KEYINPUT4), .C2(new_n436_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(new_n433_), .C1(new_n445_), .C2(new_n434_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n419_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n415_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(new_n409_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n455_), .A2(new_n458_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n452_), .A2(new_n464_), .A3(new_n432_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n452_), .B2(new_n432_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n463_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n454_), .B1(new_n468_), .B2(KEYINPUT104), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n453_), .A2(KEYINPUT33), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n462_), .B1(new_n470_), .B2(new_n465_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT104), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n382_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT27), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n455_), .A2(new_n475_), .A3(new_n461_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT106), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n455_), .A2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n422_), .A2(new_n426_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n459_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n455_), .A2(new_n477_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n476_), .B1(new_n482_), .B2(KEYINPUT27), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n376_), .A2(new_n381_), .A3(new_n377_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n451_), .A2(new_n453_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n321_), .B1(new_n474_), .B2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n382_), .A2(new_n483_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n485_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n321_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n267_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G230gat), .A2(G233gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT64), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G64gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G57gat), .ZN(new_n497_));
  INV_X1    g296(.A(G57gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G64gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT11), .ZN(new_n500_));
  INV_X1    g299(.A(G78gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G71gat), .ZN(new_n502_));
  INV_X1    g301(.A(G71gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G78gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n507_), .A2(KEYINPUT11), .A3(new_n502_), .A4(new_n504_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n245_), .A2(new_n247_), .A3(new_n511_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n495_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(KEYINPUT12), .B(new_n510_), .C1(new_n506_), .C2(new_n508_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n241_), .A2(KEYINPUT67), .A3(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(new_n514_), .C1(KEYINPUT12), .C2(new_n512_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n515_), .B1(new_n524_), .B2(new_n495_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G120gat), .B(G148gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT5), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G176gat), .B(G204gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n525_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT13), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT73), .B(G1gat), .ZN(new_n534_));
  INV_X1    g333(.A(G8gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT74), .Z(new_n539_));
  XNOR2_X1  g338(.A(G1gat), .B(G8gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n538_), .B(KEYINPUT74), .ZN(new_n542_));
  INV_X1    g341(.A(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n511_), .B(new_n546_), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n545_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT78), .Z(new_n549_));
  XOR2_X1   g348(.A(G127gat), .B(G155gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT17), .Z(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n548_), .B(KEYINPUT75), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n210_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n545_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n545_), .A2(new_n566_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n211_), .A2(new_n541_), .A3(new_n544_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n563_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n572_), .A3(new_n563_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT79), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n573_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n533_), .A2(new_n560_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n492_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n582_), .B2(new_n489_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT107), .Z(new_n584_));
  AOI21_X1  g383(.A(new_n580_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT72), .B(KEYINPUT37), .Z(new_n586_));
  NAND3_X1  g385(.A1(new_n263_), .A2(new_n265_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n259_), .A2(new_n257_), .A3(new_n255_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n206_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n264_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT70), .B1(new_n590_), .B2(KEYINPUT37), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT70), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n592_), .B(new_n593_), .C1(new_n589_), .C2(new_n264_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n587_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n596_), .A2(new_n560_), .A3(new_n533_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n585_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n485_), .A3(new_n534_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT38), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n584_), .A2(new_n601_), .ZN(G1324gat));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n535_), .A3(new_n483_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n492_), .A2(new_n483_), .A3(new_n581_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n604_), .A2(KEYINPUT108), .A3(new_n605_), .A4(G8gat), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT108), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n535_), .B1(new_n608_), .B2(KEYINPUT39), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n604_), .A2(new_n609_), .B1(KEYINPUT108), .B2(new_n605_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n603_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g411(.A(G15gat), .B1(new_n582_), .B2(new_n321_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT41), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n599_), .A2(new_n272_), .A3(new_n490_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  OAI21_X1  g415(.A(G22gat), .B1(new_n582_), .B2(new_n484_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT42), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n484_), .A2(G22gat), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n618_), .B1(new_n598_), .B2(new_n619_), .ZN(G1327gat));
  NAND2_X1  g419(.A1(new_n267_), .A2(new_n560_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n621_), .A2(new_n533_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n585_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(G29gat), .B1(new_n624_), .B2(new_n485_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT110), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n595_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n626_), .B(KEYINPUT43), .C1(new_n627_), .C2(KEYINPUT109), .ZN(new_n628_));
  INV_X1    g427(.A(new_n560_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n533_), .A2(new_n629_), .A3(new_n580_), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n471_), .A2(new_n472_), .B1(new_n489_), .B2(new_n428_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n468_), .A2(KEYINPUT104), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n484_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n480_), .A2(new_n481_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n475_), .B1(new_n634_), .B2(new_n478_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n382_), .B(new_n489_), .C1(new_n476_), .C2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n490_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n637_));
  NOR4_X1   g436(.A1(new_n382_), .A2(new_n321_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n596_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT109), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT110), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n627_), .B2(new_n626_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n628_), .B(new_n630_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT43), .B1(new_n639_), .B2(KEYINPUT110), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n626_), .B1(new_n627_), .B2(KEYINPUT109), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n628_), .A4(new_n630_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n485_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n625_), .B1(new_n652_), .B2(new_n653_), .ZN(G1328gat));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n650_), .A3(new_n483_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G36gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n483_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n623_), .A2(G36gat), .A3(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT45), .Z(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(KEYINPUT46), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  OAI21_X1  g463(.A(new_n269_), .B1(new_n623_), .B2(new_n321_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT111), .Z(new_n666_));
  NAND2_X1  g465(.A1(new_n490_), .A2(G43gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n651_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g468(.A(G50gat), .B1(new_n651_), .B2(new_n484_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n484_), .A2(G50gat), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT112), .Z(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n623_), .B2(new_n672_), .ZN(G1331gat));
  INV_X1    g472(.A(new_n580_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n596_), .A2(new_n560_), .A3(new_n532_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n489_), .B1(new_n677_), .B2(KEYINPUT113), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(KEYINPUT113), .B2(new_n677_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n674_), .A2(new_n532_), .A3(new_n560_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n492_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n498_), .B1(new_n485_), .B2(KEYINPUT114), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(KEYINPUT114), .B2(new_n498_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n679_), .A2(new_n498_), .B1(new_n682_), .B2(new_n684_), .ZN(G1332gat));
  OAI21_X1  g484(.A(G64gat), .B1(new_n681_), .B2(new_n657_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT48), .ZN(new_n687_));
  INV_X1    g486(.A(new_n677_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n496_), .A3(new_n483_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1333gat));
  OAI21_X1  g489(.A(G71gat), .B1(new_n681_), .B2(new_n321_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(new_n503_), .A3(new_n490_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1334gat));
  NAND3_X1  g494(.A1(new_n688_), .A2(new_n501_), .A3(new_n382_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n501_), .B1(new_n682_), .B2(new_n382_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT50), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n698_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT116), .Z(G1335gat));
  NOR3_X1   g502(.A1(new_n674_), .A2(new_n532_), .A3(new_n629_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT117), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n649_), .A2(new_n628_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n489_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n621_), .A2(new_n532_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n675_), .A2(new_n709_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n489_), .A2(G85gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(G1336gat));
  OAI21_X1  g511(.A(G92gat), .B1(new_n707_), .B2(new_n657_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n657_), .A2(G92gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n710_), .B2(new_n714_), .ZN(G1337gat));
  OAI21_X1  g514(.A(G99gat), .B1(new_n707_), .B2(new_n321_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n710_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n717_), .A2(new_n490_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n235_), .A3(new_n382_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n649_), .A2(new_n382_), .A3(new_n628_), .A4(new_n706_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n722_), .A2(new_n723_), .A3(G106gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n722_), .B2(G106gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n728_), .B(new_n721_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1339gat));
  NAND4_X1  g529(.A1(new_n595_), .A2(new_n629_), .A3(new_n580_), .A4(new_n532_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT54), .Z(new_n732_));
  OAI21_X1  g531(.A(new_n578_), .B1(new_n577_), .B2(new_n573_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n574_), .A2(KEYINPUT79), .A3(new_n575_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n733_), .A2(new_n734_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n518_), .A2(new_n519_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT67), .B1(new_n241_), .B2(new_n517_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n514_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n511_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT12), .B1(new_n248_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n494_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT118), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT118), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n523_), .A2(new_n743_), .A3(new_n494_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT55), .B1(new_n523_), .B2(new_n494_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n738_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n740_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .A4(new_n495_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n745_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT119), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n745_), .A2(new_n751_), .A3(KEYINPUT119), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT56), .B1(new_n756_), .B2(new_n529_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n745_), .A2(new_n751_), .A3(KEYINPUT119), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT119), .B1(new_n745_), .B2(new_n751_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT56), .B(new_n529_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n735_), .B1(new_n757_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n564_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n563_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n567_), .A2(new_n565_), .A3(new_n571_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT120), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n766_), .A2(new_n767_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n577_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n531_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n762_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n266_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT121), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n773_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT57), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT122), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n530_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(KEYINPUT56), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n529_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(KEYINPUT122), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n785_), .A3(new_n760_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n525_), .A2(new_n530_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n770_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n786_), .A2(KEYINPUT58), .A3(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n596_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT57), .B1(new_n772_), .B2(new_n266_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT121), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n777_), .A2(new_n779_), .A3(new_n793_), .A4(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n732_), .B1(new_n796_), .B2(new_n560_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n488_), .A2(new_n485_), .A3(new_n490_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT59), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n793_), .A2(new_n775_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n800_), .A2(KEYINPUT123), .B1(KEYINPUT57), .B2(new_n778_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n595_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n794_), .B1(new_n802_), .B2(new_n792_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n629_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(new_n732_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n799_), .B(new_n674_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(G113gat), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n797_), .A2(new_n798_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n674_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT124), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n810_), .A2(new_n816_), .A3(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1340gat));
  OAI21_X1  g617(.A(new_n799_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G120gat), .B1(new_n819_), .B2(new_n532_), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n532_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n811_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n821_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1341gat));
  OAI21_X1  g623(.A(G127gat), .B1(new_n819_), .B2(new_n560_), .ZN(new_n825_));
  INV_X1    g624(.A(G127gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n811_), .A2(new_n826_), .A3(new_n629_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1342gat));
  OAI21_X1  g627(.A(G134gat), .B1(new_n819_), .B2(new_n595_), .ZN(new_n829_));
  INV_X1    g628(.A(G134gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n811_), .A2(new_n830_), .A3(new_n267_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1343gat));
  NAND4_X1  g631(.A1(new_n657_), .A2(new_n485_), .A3(new_n382_), .A4(new_n321_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n797_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n674_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT125), .B(G141gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1344gat));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n533_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n629_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT61), .B(G155gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1346gat));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n834_), .A2(new_n843_), .A3(new_n267_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n797_), .A2(new_n595_), .A3(new_n833_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n843_), .ZN(G1347gat));
  INV_X1    g645(.A(G169gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n490_), .A2(new_n489_), .A3(new_n483_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n382_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n674_), .B(new_n849_), .C1(new_n806_), .C2(new_n732_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT62), .B(new_n847_), .C1(new_n850_), .C2(KEYINPUT22), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  INV_X1    g651(.A(new_n849_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n779_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n793_), .A2(new_n804_), .A3(new_n775_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n560_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n732_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n580_), .B(new_n853_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT22), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n852_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G169gat), .B1(new_n850_), .B2(KEYINPUT62), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n851_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT126), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT126), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n864_), .B(new_n851_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1348gat));
  NOR2_X1   g665(.A1(new_n807_), .A2(new_n853_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G176gat), .B1(new_n867_), .B2(new_n533_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n797_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n484_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G176gat), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n848_), .A2(new_n872_), .A3(new_n532_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n868_), .B1(new_n871_), .B2(new_n873_), .ZN(G1349gat));
  OR3_X1    g673(.A1(new_n870_), .A2(new_n560_), .A3(new_n848_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n560_), .B1(new_n285_), .B2(new_n289_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n875_), .A2(new_n284_), .B1(new_n867_), .B2(new_n876_), .ZN(G1350gat));
  NAND3_X1  g676(.A1(new_n867_), .A2(new_n392_), .A3(new_n267_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n807_), .A2(new_n595_), .A3(new_n853_), .ZN(new_n879_));
  INV_X1    g678(.A(G190gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(G1351gat));
  XOR2_X1   g680(.A(KEYINPUT127), .B(G197gat), .Z(new_n882_));
  NOR2_X1   g681(.A1(KEYINPUT127), .A2(G197gat), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n490_), .A2(new_n657_), .A3(new_n485_), .A4(new_n484_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n869_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n580_), .ZN(new_n886_));
  MUX2_X1   g685(.A(new_n882_), .B(new_n883_), .S(new_n886_), .Z(G1352gat));
  INV_X1    g686(.A(new_n885_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n533_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n629_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  AND2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n891_), .B2(new_n892_), .ZN(G1354gat));
  OR3_X1    g694(.A1(new_n885_), .A2(G218gat), .A3(new_n266_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G218gat), .B1(new_n885_), .B2(new_n595_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1355gat));
endmodule


