//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_;
  XNOR2_X1  g000(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  AND2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT72), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G29gat), .ZN(new_n207_));
  INV_X1    g006(.A(G36gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G43gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n206_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n206_), .B2(new_n212_), .ZN(new_n215_));
  INV_X1    g014(.A(G50gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT72), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n210_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n219_));
  OAI21_X1  g018(.A(G43gat), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n206_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n221_));
  AOI21_X1  g020(.A(G50gat), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n203_), .B1(new_n217_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n216_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(G50gat), .A3(new_n221_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n202_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(G15gat), .ZN(new_n228_));
  INV_X1    g027(.A(G22gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G1gat), .ZN(new_n231_));
  INV_X1    g030(.A(G8gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT14), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G1gat), .B(G8gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n234_), .B(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n227_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT84), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n217_), .A2(new_n222_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT85), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n234_), .B(new_n235_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n241_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G229gat), .A3(G233gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n245_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n246_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253_));
  INV_X1    g052(.A(G169gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n252_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT65), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT7), .ZN(new_n271_));
  INV_X1    g070(.A(G99gat), .ZN(new_n272_));
  INV_X1    g071(.A(G106gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n262_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n270_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G85gat), .A2(G92gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT8), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n274_), .A2(new_n268_), .A3(new_n269_), .A4(new_n262_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n279_), .A2(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n281_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT9), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n278_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n279_), .A2(KEYINPUT9), .ZN(new_n292_));
  INV_X1    g091(.A(new_n280_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n278_), .A2(KEYINPUT64), .A3(new_n288_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT10), .B(G99gat), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n273_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n270_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n283_), .A2(new_n287_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT66), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n277_), .A2(new_n282_), .B1(new_n286_), .B2(new_n281_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G57gat), .B(G64gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT11), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G71gat), .B(G78gat), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n305_), .A2(KEYINPUT11), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n307_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n304_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT67), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(KEYINPUT67), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G230gat), .A2(G233gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n261_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n314_), .A2(KEYINPUT67), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n314_), .A2(KEYINPUT67), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT68), .B(new_n320_), .C1(new_n323_), .C2(new_n313_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n283_), .A2(new_n326_), .A3(new_n287_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n298_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n311_), .B(KEYINPUT70), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT12), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n313_), .B2(KEYINPUT12), .ZN(new_n332_));
  OR3_X1    g131(.A1(new_n332_), .A2(new_n314_), .A3(new_n320_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G120gat), .B(G148gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT5), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G176gat), .ZN(new_n337_));
  INV_X1    g136(.A(G204gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n325_), .A2(new_n333_), .A3(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(KEYINPUT71), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n325_), .B2(new_n333_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n332_), .A2(new_n314_), .A3(new_n320_), .ZN(new_n346_));
  AOI211_X1 g145(.A(new_n346_), .B(new_n339_), .C1(new_n319_), .C2(new_n324_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n344_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT13), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n343_), .A2(new_n348_), .A3(KEYINPUT13), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n260_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354_));
  INV_X1    g153(.A(G141gat), .ZN(new_n355_));
  INV_X1    g154(.A(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT1), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n354_), .B(new_n357_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n363_), .A2(new_n355_), .A3(new_n356_), .A4(KEYINPUT89), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT89), .ZN(new_n365_));
  OAI22_X1  g164(.A1(new_n365_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n354_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n362_), .B(new_n358_), .C1(new_n367_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n361_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G120gat), .ZN(new_n374_));
  INV_X1    g173(.A(G113gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G127gat), .A2(G134gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G127gat), .A2(G134gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n380_), .A2(new_n376_), .A3(G113gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n374_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n375_), .A3(new_n378_), .ZN(new_n383_));
  OAI21_X1  g182(.A(G113gat), .B1(new_n380_), .B2(new_n376_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(G120gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n373_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT100), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n361_), .A2(new_n382_), .A3(new_n372_), .A4(new_n385_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n386_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n391_), .A2(KEYINPUT100), .A3(new_n372_), .A4(new_n361_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT101), .B1(new_n387_), .B2(KEYINPUT4), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n387_), .A2(KEYINPUT101), .A3(KEYINPUT4), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n396_), .B(new_n398_), .C1(new_n393_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n394_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n395_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT103), .B(G1gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(new_n207_), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n405_), .B(new_n407_), .Z(new_n408_));
  NAND2_X1  g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n393_), .A2(new_n394_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n399_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n396_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n397_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n410_), .B1(new_n413_), .B2(new_n394_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n408_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(G64gat), .ZN(new_n420_));
  INV_X1    g219(.A(G92gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT104), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n425_));
  XOR2_X1   g224(.A(G211gat), .B(G218gat), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G197gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n338_), .A2(G197gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n427_), .B1(new_n434_), .B2(KEYINPUT93), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT21), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n432_), .B1(new_n430_), .B2(G197gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT93), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n426_), .B1(new_n437_), .B2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n430_), .A2(new_n256_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G197gat), .A2(G204gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(KEYINPUT21), .A3(new_n442_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n435_), .A2(new_n439_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT96), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT96), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT26), .B(G190gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n451_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT23), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT23), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(G183gat), .A3(G190gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  MUX2_X1   g264(.A(new_n465_), .B(new_n464_), .S(KEYINPUT86), .Z(new_n466_));
  NOR2_X1   g265(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G169gat), .ZN(new_n468_));
  INV_X1    g267(.A(G183gat), .ZN(new_n469_));
  INV_X1    g268(.A(G190gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n460_), .A2(new_n466_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n425_), .B1(new_n444_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n463_), .A2(KEYINPUT86), .A3(G183gat), .A4(G190gat), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n471_), .B(new_n476_), .C1(new_n465_), .C2(KEYINPUT86), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n468_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n449_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n454_), .A2(new_n459_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n465_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n475_), .B1(new_n444_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n458_), .A2(new_n459_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n466_), .A3(new_n479_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n472_), .A2(new_n468_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n437_), .A2(new_n438_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n256_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT93), .B1(new_n490_), .B2(new_n432_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n489_), .A2(KEYINPUT21), .A3(new_n426_), .A4(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n431_), .A2(new_n436_), .A3(new_n433_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n443_), .A2(new_n493_), .A3(new_n427_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(KEYINPUT97), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G226gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT19), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n474_), .A2(new_n484_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n482_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n486_), .A2(new_n492_), .A3(new_n494_), .A4(new_n487_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT20), .ZN(new_n502_));
  INV_X1    g301(.A(new_n498_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n423_), .A2(KEYINPUT104), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n424_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n474_), .A2(new_n484_), .A3(new_n496_), .A4(new_n503_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n502_), .A2(new_n498_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n423_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n417_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT98), .B1(new_n505_), .B2(new_n422_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n505_), .A2(new_n422_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n422_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT98), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n515_), .A2(new_n499_), .A3(new_n504_), .A4(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n513_), .A2(KEYINPUT99), .A3(new_n514_), .A4(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n415_), .B1(new_n413_), .B2(new_n394_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n394_), .B2(new_n393_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n402_), .A2(KEYINPUT33), .A3(new_n408_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT33), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n512_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n530_));
  XOR2_X1   g329(.A(G22gat), .B(G50gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n530_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(G228gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(G228gat), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n535_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n495_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n373_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n495_), .B2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G78gat), .B(G106gat), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n543_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n534_), .B1(new_n549_), .B2(KEYINPUT95), .ZN(new_n550_));
  INV_X1    g349(.A(new_n546_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n495_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n548_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT95), .A4(new_n534_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G227gat), .A2(G233gat), .ZN(new_n560_));
  INV_X1    g359(.A(G15gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G43gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G71gat), .B(G99gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT30), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n478_), .A2(new_n481_), .A3(new_n565_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n563_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n563_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n566_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT87), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n570_), .B2(new_n566_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT87), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n386_), .B(KEYINPUT31), .Z(new_n578_));
  AND3_X1   g377(.A1(new_n573_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n573_), .A2(new_n578_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT88), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n573_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n582_), .B(new_n583_), .C1(new_n573_), .C2(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n559_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n529_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n558_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n579_), .A2(new_n580_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n557_), .A3(new_n556_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n510_), .A2(new_n515_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n514_), .A2(new_n592_), .A3(KEYINPUT27), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT27), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(new_n518_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n417_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n591_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n587_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n353_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n601_));
  INV_X1    g400(.A(new_n298_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n283_), .A2(new_n287_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT69), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n301_), .A2(new_n326_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n601_), .B1(new_n606_), .B2(new_n227_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n224_), .A2(new_n225_), .A3(new_n202_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n202_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n329_), .A3(KEYINPUT74), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT76), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n241_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n614_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n613_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n613_), .B1(new_n612_), .B2(new_n619_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(G134gat), .ZN(new_n626_));
  INV_X1    g425(.A(G162gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT75), .B1(new_n614_), .B2(new_n618_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n299_), .A2(KEYINPUT66), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n302_), .B1(new_n301_), .B2(new_n298_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n242_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT75), .ZN(new_n633_));
  INV_X1    g432(.A(new_n618_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n606_), .A2(new_n227_), .A3(new_n601_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT74), .B1(new_n610_), .B2(new_n329_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n629_), .B(new_n635_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n617_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n623_), .A2(new_n624_), .A3(new_n628_), .A4(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n619_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT76), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n642_), .A3(new_n620_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n628_), .A2(new_n624_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n628_), .A2(new_n624_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n247_), .B(new_n311_), .ZN(new_n648_));
  AND2_X1   g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n649_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT70), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G127gat), .B(G155gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT16), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(new_n469_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(G211gat), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT17), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT70), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n650_), .A2(new_n660_), .A3(new_n651_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n653_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT80), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT82), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n652_), .A2(KEYINPUT81), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT81), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n650_), .A2(new_n666_), .A3(new_n651_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n657_), .B(new_n658_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n664_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT82), .B(new_n669_), .C1(new_n665_), .C2(new_n667_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n663_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n600_), .A2(new_n647_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n596_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT83), .B1(new_n663_), .B2(new_n673_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT80), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n662_), .B(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT83), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n679_), .B(new_n680_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n677_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n644_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT78), .Z(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n647_), .A2(new_n684_), .A3(new_n689_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n599_), .A2(new_n682_), .A3(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n695_), .A2(new_n231_), .A3(new_n417_), .A4(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT38), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n676_), .B1(new_n701_), .B2(new_n702_), .ZN(G1324gat));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n675_), .B2(new_n595_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n647_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n674_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n599_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n595_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(KEYINPUT107), .A3(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n705_), .A2(G8gat), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT39), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT39), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n705_), .A2(new_n713_), .A3(G8gat), .A4(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n695_), .A2(new_n696_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n232_), .A3(new_n709_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT40), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(KEYINPUT40), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1325gat));
  INV_X1    g521(.A(new_n581_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n584_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n716_), .A2(new_n561_), .A3(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT108), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n561_), .B1(new_n708_), .B2(new_n726_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT41), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1326gat));
  NAND3_X1  g530(.A1(new_n716_), .A2(new_n229_), .A3(new_n558_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G22gat), .B1(new_n675_), .B2(new_n559_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT42), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1327gat));
  NAND2_X1  g534(.A1(new_n682_), .A2(new_n706_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n599_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n207_), .A3(new_n417_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n691_), .A2(new_n692_), .B1(new_n587_), .B2(new_n597_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n739_), .B2(KEYINPUT109), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n689_), .B1(new_n647_), .B2(new_n684_), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n683_), .B(new_n690_), .C1(new_n640_), .C2(new_n646_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT33), .B1(new_n402_), .B2(new_n408_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n414_), .A2(new_n526_), .A3(new_n415_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n745_), .A2(new_n520_), .A3(new_n524_), .A4(new_n521_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n585_), .B1(new_n746_), .B2(new_n512_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n591_), .A2(new_n596_), .A3(new_n595_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n741_), .A2(new_n742_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n740_), .A2(new_n353_), .A3(new_n682_), .A4(new_n752_), .ZN(new_n753_));
  OR2_X1    g552(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n754_));
  NAND2_X1  g553(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT111), .B1(new_n753_), .B2(new_n758_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n751_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n677_), .A2(new_n681_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(KEYINPUT44), .A4(new_n353_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n757_), .B1(new_n759_), .B2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(new_n417_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n738_), .B1(new_n767_), .B2(new_n207_), .ZN(G1328gat));
  NAND3_X1  g567(.A1(new_n737_), .A2(new_n208_), .A3(new_n709_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT45), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n756_), .A2(new_n709_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n765_), .A2(new_n759_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n774_), .B2(G36gat), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT112), .B(new_n208_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n770_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n770_), .B(KEYINPUT46), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1329gat));
  INV_X1    g580(.A(new_n737_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n213_), .B1(new_n782_), .B2(new_n725_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n579_), .A2(new_n213_), .A3(new_n580_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT113), .B1(new_n766_), .B2(new_n784_), .ZN(new_n785_));
  AND4_X1   g584(.A1(KEYINPUT113), .A2(new_n773_), .A3(new_n756_), .A4(new_n784_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT47), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n789_), .B(new_n783_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1330gat));
  NAND3_X1  g590(.A1(new_n737_), .A2(new_n216_), .A3(new_n558_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n766_), .A2(new_n558_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n216_), .ZN(G1331gat));
  AND3_X1   g593(.A1(new_n343_), .A2(new_n348_), .A3(KEYINPUT13), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT13), .B1(new_n343_), .B2(new_n348_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n259_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n598_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n798_), .A2(new_n682_), .A3(new_n693_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G57gat), .B1(new_n799_), .B2(new_n417_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(KEYINPUT114), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(KEYINPUT114), .ZN(new_n802_));
  INV_X1    g601(.A(new_n798_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n647_), .A3(new_n762_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n417_), .A2(G57gat), .ZN(new_n805_));
  OAI22_X1  g604(.A1(new_n801_), .A2(new_n802_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT115), .Z(G1332gat));
  OAI21_X1  g606(.A(G64gat), .B1(new_n804_), .B2(new_n595_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT48), .ZN(new_n809_));
  INV_X1    g608(.A(G64gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n799_), .A2(new_n810_), .A3(new_n709_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1333gat));
  OAI21_X1  g611(.A(G71gat), .B1(new_n804_), .B2(new_n725_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT49), .ZN(new_n816_));
  INV_X1    g615(.A(G71gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n799_), .A2(new_n817_), .A3(new_n726_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1334gat));
  OAI21_X1  g618(.A(G78gat), .B1(new_n804_), .B2(new_n559_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G78gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n799_), .A2(new_n823_), .A3(new_n558_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1335gat));
  NOR2_X1   g624(.A1(new_n798_), .A2(new_n736_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G85gat), .B1(new_n826_), .B2(new_n417_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n740_), .A2(new_n682_), .A3(new_n797_), .A4(new_n752_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT118), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n417_), .A2(G85gat), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT119), .Z(new_n835_));
  AOI21_X1  g634(.A(new_n827_), .B1(new_n833_), .B2(new_n835_), .ZN(G1336gat));
  AOI21_X1  g635(.A(G92gat), .B1(new_n826_), .B2(new_n709_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n595_), .A2(new_n421_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n833_), .B2(new_n838_), .ZN(G1337gat));
  NAND3_X1  g638(.A1(new_n830_), .A2(new_n726_), .A3(new_n832_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G99gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n589_), .A2(new_n296_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n826_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n841_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT121), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n841_), .A2(new_n850_), .A3(new_n847_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT51), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n841_), .B2(new_n847_), .ZN(new_n853_));
  AOI211_X1 g652(.A(KEYINPUT121), .B(new_n846_), .C1(new_n840_), .C2(G99gat), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n852_), .A2(new_n856_), .ZN(G1338gat));
  NAND3_X1  g656(.A1(new_n826_), .A2(new_n273_), .A3(new_n558_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n829_), .A2(new_n558_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(G106gat), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n859_), .B2(G106gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n858_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n333_), .B2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n346_), .A2(KEYINPUT122), .A3(KEYINPUT55), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n320_), .B1(new_n323_), .B2(new_n332_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n346_), .B1(new_n872_), .B2(KEYINPUT55), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n339_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT56), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n339_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n259_), .A2(new_n875_), .A3(new_n342_), .A4(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n249_), .A2(new_n240_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n239_), .A2(new_n243_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n240_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n258_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n252_), .B2(new_n258_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n343_), .A2(new_n348_), .A3(new_n883_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n878_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT123), .B(new_n866_), .C1(new_n885_), .C2(new_n706_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n875_), .A2(new_n877_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n342_), .A3(new_n883_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n887_), .A2(KEYINPUT58), .A3(new_n342_), .A4(new_n883_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n693_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n706_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(KEYINPUT57), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(KEYINPUT57), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n886_), .A2(new_n892_), .A3(new_n895_), .A4(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n707_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n682_), .A2(new_n693_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n795_), .A2(new_n796_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n260_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT54), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n899_), .A2(new_n904_), .A3(new_n260_), .A4(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n898_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n709_), .A2(new_n596_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n590_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n907_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G113gat), .B1(new_n913_), .B2(new_n259_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(KEYINPUT59), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n892_), .A2(new_n896_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n894_), .A2(KEYINPUT57), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n682_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n906_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n919_), .A2(new_n920_), .A3(new_n911_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n915_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n260_), .A2(new_n375_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n914_), .B1(new_n922_), .B2(new_n923_), .ZN(G1340gat));
  NAND3_X1  g723(.A1(new_n915_), .A2(new_n900_), .A3(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(G120gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n374_), .B1(new_n901_), .B2(KEYINPUT60), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n913_), .B(new_n927_), .C1(KEYINPUT60), .C2(new_n374_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1341gat));
  AOI21_X1  g728(.A(G127gat), .B1(new_n913_), .B2(new_n762_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n674_), .A2(G127gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n922_), .B2(new_n931_), .ZN(G1342gat));
  AOI21_X1  g731(.A(G134gat), .B1(new_n913_), .B2(new_n706_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n693_), .A2(G134gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n922_), .B2(new_n934_), .ZN(G1343gat));
  INV_X1    g734(.A(new_n588_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n907_), .A2(new_n936_), .A3(new_n908_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n259_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(G141gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n937_), .A2(new_n355_), .A3(new_n259_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1344gat));
  NAND2_X1  g740(.A1(new_n937_), .A2(new_n900_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(G148gat), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n937_), .A2(new_n356_), .A3(new_n900_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1345gat));
  NAND4_X1  g744(.A1(new_n907_), .A2(new_n936_), .A3(new_n762_), .A4(new_n908_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT61), .B(G155gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n946_), .B(new_n947_), .ZN(G1346gat));
  AOI21_X1  g747(.A(G162gat), .B1(new_n937_), .B2(new_n706_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n693_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(new_n627_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n937_), .B2(new_n951_), .ZN(G1347gat));
  NOR4_X1   g751(.A1(new_n595_), .A2(new_n725_), .A3(new_n417_), .A4(new_n558_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n918_), .B2(new_n906_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT22), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n955_), .A2(new_n956_), .A3(new_n259_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n957_), .A2(KEYINPUT62), .A3(new_n254_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n919_), .A2(new_n953_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n959_), .A2(KEYINPUT62), .A3(new_n260_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n960_), .A2(new_n254_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n957_), .A2(KEYINPUT62), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n958_), .B1(new_n961_), .B2(new_n962_), .ZN(G1348gat));
  AOI21_X1  g762(.A(G176gat), .B1(new_n955_), .B2(new_n900_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n897_), .A2(new_n707_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n965_), .A2(new_n954_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n900_), .A2(G176gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n964_), .B1(new_n966_), .B2(new_n967_), .ZN(G1349gat));
  NOR3_X1   g767(.A1(new_n959_), .A2(new_n458_), .A3(new_n707_), .ZN(new_n969_));
  AOI21_X1  g768(.A(KEYINPUT124), .B1(new_n966_), .B2(new_n762_), .ZN(new_n970_));
  AND4_X1   g769(.A1(KEYINPUT124), .A2(new_n907_), .A3(new_n762_), .A4(new_n953_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n969_), .B1(new_n972_), .B2(new_n469_), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n955_), .A2(new_n706_), .A3(new_n459_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n955_), .A2(new_n693_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n975_), .B1(new_n976_), .B2(G190gat), .ZN(new_n977_));
  AOI211_X1 g776(.A(KEYINPUT125), .B(new_n470_), .C1(new_n955_), .C2(new_n693_), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n974_), .B1(new_n977_), .B2(new_n978_), .ZN(G1351gat));
  NAND2_X1  g778(.A1(new_n936_), .A2(new_n596_), .ZN(new_n980_));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n980_), .A2(new_n981_), .ZN(new_n982_));
  NOR2_X1   g781(.A1(new_n965_), .A2(new_n982_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n595_), .B1(new_n980_), .B2(new_n981_), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n983_), .A2(new_n259_), .A3(new_n984_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g785(.A(new_n982_), .ZN(new_n987_));
  AND3_X1   g786(.A1(new_n907_), .A2(new_n987_), .A3(new_n984_), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n988_), .A2(new_n900_), .A3(new_n430_), .ZN(new_n989_));
  AND2_X1   g788(.A1(new_n988_), .A2(new_n900_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n990_), .B2(new_n338_), .ZN(G1353gat));
  NAND2_X1  g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  NAND4_X1  g791(.A1(new_n983_), .A2(new_n674_), .A3(new_n984_), .A4(new_n992_), .ZN(new_n993_));
  NOR2_X1   g792(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n994_));
  XNOR2_X1  g793(.A(new_n994_), .B(KEYINPUT127), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n993_), .B(new_n995_), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n988_), .B2(new_n706_), .ZN(new_n997_));
  AND2_X1   g796(.A1(new_n693_), .A2(G218gat), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n997_), .B1(new_n988_), .B2(new_n998_), .ZN(G1355gat));
endmodule


