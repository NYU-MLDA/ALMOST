//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_;
  INV_X1    g000(.A(KEYINPUT26), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT95), .B1(new_n203_), .B2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n202_), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT95), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n207_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT96), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(KEYINPUT96), .A3(KEYINPUT24), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n222_), .B1(new_n223_), .B2(new_n204_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n212_), .A2(new_n221_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT97), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n212_), .A2(new_n228_), .A3(KEYINPUT97), .A4(new_n221_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G204gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT90), .B1(new_n234_), .B2(G197gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236_));
  INV_X1    g035(.A(G197gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(G204gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT21), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(G197gat), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .A4(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n234_), .A2(G197gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n237_), .A2(G204gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT21), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G218gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G211gat), .ZN(new_n246_));
  INV_X1    g045(.A(G211gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G218gat), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT91), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT91), .B1(new_n246_), .B2(new_n248_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n241_), .B(new_n244_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n248_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT91), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n235_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT91), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT21), .A4(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n251_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n223_), .A2(new_n204_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n224_), .A2(new_n259_), .A3(new_n225_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n213_), .A2(KEYINPUT83), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(G169gat), .A3(G176gat), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(KEYINPUT84), .A2(G176gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n217_), .A2(KEYINPUT22), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT22), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(KEYINPUT84), .A2(G176gat), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n265_), .A2(new_n266_), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n264_), .A2(new_n270_), .A3(KEYINPUT98), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT98), .B1(new_n264_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n260_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n233_), .A2(new_n258_), .A3(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n207_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT82), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n261_), .A2(new_n263_), .A3(new_n219_), .A4(KEYINPUT24), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT82), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n207_), .A2(new_n280_), .A3(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n282_), .A2(new_n228_), .A3(new_n283_), .A4(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n270_), .A2(KEYINPUT85), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT85), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT84), .A2(G176gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT84), .A2(G176gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G169gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n288_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n264_), .B1(new_n287_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n260_), .A2(KEYINPUT86), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT86), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n224_), .A2(new_n259_), .A3(new_n296_), .A4(new_n225_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n286_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n251_), .A2(new_n257_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n279_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n274_), .A2(new_n278_), .A3(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G8gat), .B(G36gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n270_), .A2(KEYINPUT85), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n291_), .A2(new_n292_), .A3(new_n288_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n312_), .A2(new_n264_), .A3(new_n295_), .A4(new_n297_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n258_), .A2(new_n313_), .A3(new_n286_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT20), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n233_), .A2(new_n273_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n300_), .ZN(new_n319_));
  OAI211_X1 g118(.A(KEYINPUT94), .B(KEYINPUT20), .C1(new_n299_), .C2(new_n300_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n321_), .A2(KEYINPUT99), .A3(new_n277_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT99), .B1(new_n321_), .B2(new_n277_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n302_), .B(new_n309_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n258_), .A2(new_n273_), .A3(new_n229_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n301_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n277_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n321_), .B2(new_n277_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n309_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  OR2_X1    g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G141gat), .ZN(new_n338_));
  INV_X1    g137(.A(G148gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT88), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n338_), .B(new_n339_), .C1(new_n340_), .C2(KEYINPUT3), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n342_), .B(KEYINPUT88), .C1(G141gat), .C2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n341_), .A2(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n349_), .A2(KEYINPUT2), .B1(new_n340_), .B2(KEYINPUT3), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n337_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT87), .B1(new_n336_), .B2(KEYINPUT1), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(G155gat), .A4(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n336_), .A2(KEYINPUT1), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n352_), .A2(new_n355_), .A3(new_n335_), .A4(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G141gat), .B(G148gat), .Z(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n334_), .B1(new_n351_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n341_), .A2(new_n343_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n345_), .A2(new_n344_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n350_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n337_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n357_), .A2(new_n358_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n332_), .B(new_n333_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n368_), .A3(KEYINPUT101), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n351_), .A2(new_n359_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT101), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(KEYINPUT4), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n360_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT102), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n369_), .A2(new_n372_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT103), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n380_), .A2(KEYINPUT103), .A3(new_n381_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n379_), .A2(new_n384_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT103), .B1(new_n380_), .B2(new_n381_), .ZN(new_n392_));
  AOI211_X1 g191(.A(new_n383_), .B(new_n378_), .C1(new_n369_), .C2(new_n372_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n388_), .B1(new_n394_), .B2(new_n379_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n331_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT106), .B1(new_n325_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n379_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n388_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n400_), .A2(new_n390_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT106), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n324_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n302_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n307_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n380_), .A2(KEYINPUT104), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT104), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n369_), .A2(new_n408_), .A3(new_n372_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n381_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n378_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n410_), .A2(new_n388_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n390_), .A2(KEYINPUT33), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n394_), .A2(new_n414_), .A3(new_n388_), .A4(new_n379_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n308_), .B(new_n302_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n406_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT105), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT105), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n406_), .A2(new_n416_), .A3(new_n420_), .A4(new_n417_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n404_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n300_), .B1(new_n370_), .B2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(G228gat), .A2(G233gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(KEYINPUT92), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G78gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G106gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n428_), .B(G78gat), .ZN(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n424_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n370_), .A2(new_n425_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT28), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n427_), .A2(KEYINPUT92), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n431_), .A2(new_n434_), .A3(new_n424_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n440_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n435_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT107), .B1(new_n422_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n400_), .A2(new_n390_), .ZN(new_n449_));
  AND4_X1   g248(.A1(new_n402_), .A2(new_n324_), .A3(new_n449_), .A4(new_n331_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n402_), .B1(new_n401_), .B2(new_n324_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT99), .ZN(new_n453_));
  INV_X1    g252(.A(new_n320_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT94), .B1(new_n314_), .B2(KEYINPUT20), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n258_), .B1(new_n233_), .B2(new_n273_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n453_), .B1(new_n457_), .B2(new_n278_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n321_), .A2(KEYINPUT99), .A3(new_n277_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n308_), .B1(new_n460_), .B2(new_n302_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n302_), .ZN(new_n462_));
  AOI211_X1 g261(.A(new_n307_), .B(new_n462_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n420_), .B1(new_n464_), .B2(new_n416_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n421_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n452_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT107), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n446_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n449_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n461_), .A2(new_n463_), .A3(KEYINPUT27), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n329_), .A2(new_n307_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT108), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n417_), .B2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n460_), .A2(KEYINPUT108), .A3(new_n308_), .A4(new_n302_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n447_), .B(new_n470_), .C1(new_n471_), .C2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n448_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G43gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n299_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(new_n367_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(G15gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT30), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT31), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n483_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n446_), .B1(new_n477_), .B2(new_n471_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT109), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT109), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n446_), .B(new_n493_), .C1(new_n477_), .C2(new_n471_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n492_), .A2(new_n494_), .A3(new_n489_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n479_), .A2(new_n490_), .B1(new_n495_), .B2(new_n470_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497_));
  INV_X1    g296(.A(G1gat), .ZN(new_n498_));
  INV_X1    g297(.A(G8gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n497_), .B1(new_n500_), .B2(KEYINPUT75), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n500_), .A2(KEYINPUT75), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G1gat), .B(G8gat), .ZN(new_n503_));
  OR3_X1    g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G29gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(KEYINPUT15), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n505_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT80), .Z(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n511_), .B(new_n508_), .Z(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(G229gat), .A3(G233gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT79), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n515_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n518_), .B2(new_n517_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G113gat), .B(G141gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT81), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G169gat), .B(G197gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n520_), .B(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT6), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n528_));
  OR3_X1    g327(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G85gat), .B(G92gat), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT64), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT64), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n530_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT8), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(KEYINPUT9), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT10), .B(G99gat), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n433_), .ZN(new_n540_));
  INV_X1    g339(.A(G85gat), .ZN(new_n541_));
  INV_X1    g340(.A(G92gat), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n541_), .A2(new_n542_), .A3(KEYINPUT9), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(new_n540_), .A3(new_n527_), .A4(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n537_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G57gat), .B(G64gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT11), .ZN(new_n547_));
  XOR2_X1   g346(.A(G71gat), .B(G78gat), .Z(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n546_), .A2(KEYINPUT11), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n548_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n545_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT12), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n545_), .A2(new_n552_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n545_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n555_), .A2(KEYINPUT65), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n553_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n545_), .A2(KEYINPUT65), .A3(new_n552_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n563_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G120gat), .B(G148gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n561_), .A2(new_n565_), .A3(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(KEYINPUT67), .Z(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT13), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT68), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(KEYINPUT68), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n571_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n496_), .A2(new_n525_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n545_), .A2(new_n508_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT34), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n537_), .A2(new_n544_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n588_), .A2(KEYINPUT70), .A3(new_n510_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT70), .B1(new_n588_), .B2(new_n510_), .ZN(new_n590_));
  OAI221_X1 g389(.A(new_n585_), .B1(KEYINPUT35), .B2(new_n587_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(KEYINPUT35), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT69), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n591_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n593_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n591_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT74), .ZN(new_n599_));
  XOR2_X1   g398(.A(G190gat), .B(G218gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT71), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT73), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n599_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n604_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT72), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n594_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n598_), .A2(new_n606_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n614_), .A3(KEYINPUT37), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n552_), .B(new_n617_), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT76), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n511_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n620_), .A2(KEYINPUT78), .ZN(new_n627_));
  INV_X1    g426(.A(new_n625_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n626_), .A2(KEYINPUT17), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n627_), .A2(KEYINPUT17), .A3(new_n628_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n616_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n584_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n498_), .A3(new_n449_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT38), .ZN(new_n635_));
  INV_X1    g434(.A(new_n611_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n631_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n584_), .A2(KEYINPUT110), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n419_), .A2(new_n421_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n447_), .B1(new_n639_), .B2(new_n452_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n478_), .B1(new_n640_), .B2(new_n468_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n422_), .A2(KEYINPUT107), .A3(new_n447_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n490_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n495_), .A2(new_n470_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n583_), .A2(new_n525_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n637_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT110), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n470_), .B1(new_n638_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n635_), .B1(new_n650_), .B2(new_n498_), .ZN(G1324gat));
  NOR2_X1   g450(.A1(new_n477_), .A2(new_n471_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n633_), .A2(new_n499_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G8gat), .B1(new_n647_), .B2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g458(.A1(new_n638_), .A2(new_n649_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n489_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT111), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(G15gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n490_), .B1(new_n638_), .B2(new_n649_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT111), .B1(new_n664_), .B2(new_n485_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(KEYINPUT41), .A3(new_n665_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n633_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT112), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n669_), .A3(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n633_), .A2(new_n673_), .A3(new_n447_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n446_), .B1(new_n638_), .B2(new_n649_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(new_n673_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT42), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT42), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1327gat));
  INV_X1    g478(.A(new_n631_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n611_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n584_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n449_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n616_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n496_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n442_), .A2(new_n445_), .A3(new_n470_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n652_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n467_), .A2(new_n446_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(KEYINPUT107), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n489_), .B1(new_n690_), .B2(new_n469_), .ZN(new_n691_));
  AND4_X1   g490(.A1(new_n470_), .A2(new_n492_), .A3(new_n494_), .A4(new_n489_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n686_), .B(new_n616_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n685_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n646_), .A2(new_n631_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n698_), .B(new_n695_), .C1(new_n685_), .C2(new_n693_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n449_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n683_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n584_), .A2(new_n703_), .A3(new_n652_), .A4(new_n681_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n697_), .A2(new_n699_), .A3(new_n654_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n703_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n705_), .B(new_n708_), .C1(new_n706_), .C2(new_n703_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  AOI21_X1  g511(.A(G43gat), .B1(new_n682_), .B2(new_n489_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n489_), .A2(G43gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n700_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1330gat));
  INV_X1    g516(.A(G50gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n682_), .A2(new_n718_), .A3(new_n447_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n700_), .A2(new_n720_), .A3(new_n447_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n700_), .B2(new_n447_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1331gat));
  INV_X1    g523(.A(new_n525_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n496_), .A2(new_n725_), .A3(new_n582_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n632_), .ZN(new_n727_));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n449_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n726_), .A2(new_n637_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n449_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n731_), .B2(new_n728_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n730_), .B2(new_n652_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT48), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n727_), .A2(new_n733_), .A3(new_n652_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n730_), .B2(new_n489_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT49), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n727_), .A2(new_n738_), .A3(new_n489_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1334gat));
  AOI21_X1  g541(.A(new_n429_), .B1(new_n730_), .B2(new_n447_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT50), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n727_), .A2(new_n429_), .A3(new_n447_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n582_), .A2(new_n725_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n631_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n694_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n470_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n726_), .A2(new_n681_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n541_), .A3(new_n449_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1336gat));
  OAI21_X1  g553(.A(G92gat), .B1(new_n750_), .B2(new_n654_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n542_), .A3(new_n652_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n752_), .A2(new_n539_), .A3(new_n489_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n750_), .A2(new_n490_), .ZN(new_n759_));
  INV_X1    g558(.A(G99gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g561(.A(new_n686_), .B1(new_n645_), .B2(new_n616_), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT43), .B(new_n684_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n447_), .B(new_n749_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n694_), .A2(KEYINPUT116), .A3(new_n447_), .A4(new_n749_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n767_), .A2(KEYINPUT52), .A3(new_n768_), .A4(G106gat), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n726_), .A2(new_n433_), .A3(new_n447_), .A4(new_n681_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n446_), .B(new_n748_), .C1(new_n685_), .C2(new_n693_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n433_), .B1(new_n774_), .B2(KEYINPUT116), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(new_n775_), .B2(new_n767_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT53), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  INV_X1    g577(.A(new_n767_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n768_), .A2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n769_), .A4(new_n772_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n783_), .ZN(G1339gat));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  INV_X1    g584(.A(new_n524_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n516_), .A2(new_n514_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n514_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n512_), .B2(new_n788_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n520_), .A2(new_n786_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n574_), .A2(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n556_), .A2(new_n557_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT118), .B1(new_n792_), .B2(new_n559_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n559_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n558_), .A2(new_n795_), .A3(new_n560_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n793_), .A2(new_n794_), .A3(new_n796_), .A4(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n799_), .A2(new_n572_), .B1(KEYINPUT119), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n725_), .A2(new_n571_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n572_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(KEYINPUT119), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n791_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n785_), .B1(new_n807_), .B2(new_n636_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(new_n809_), .A3(KEYINPUT56), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n800_), .A2(KEYINPUT120), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n799_), .A2(new_n572_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n571_), .A2(new_n790_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n810_), .A2(KEYINPUT58), .A3(new_n813_), .A4(new_n814_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n616_), .A3(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n804_), .A2(new_n805_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n820_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT57), .B(new_n611_), .C1(new_n821_), .C2(new_n791_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n808_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n631_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n631_), .A2(new_n725_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n825_), .A2(new_n826_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n631_), .B2(new_n725_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT54), .B1(new_n829_), .B2(new_n616_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n684_), .A2(new_n827_), .A3(new_n831_), .A4(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n824_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n449_), .A3(new_n495_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836_), .B2(new_n525_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n835_), .B(KEYINPUT121), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n725_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n836_), .B2(new_n582_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n582_), .A2(KEYINPUT60), .ZN(new_n843_));
  MUX2_X1   g642(.A(new_n843_), .B(KEYINPUT60), .S(G120gat), .Z(new_n844_));
  NAND2_X1  g643(.A1(new_n838_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n842_), .A2(new_n845_), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n836_), .B2(new_n631_), .ZN(new_n847_));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n838_), .A2(new_n848_), .A3(new_n680_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1342gat));
  NAND2_X1  g649(.A1(new_n838_), .A2(new_n636_), .ZN(new_n851_));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  INV_X1    g651(.A(new_n836_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n616_), .A2(G134gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT122), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n851_), .A2(new_n852_), .B1(new_n853_), .B2(new_n855_), .ZN(G1343gat));
  NAND2_X1  g655(.A1(new_n447_), .A2(new_n490_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n652_), .A3(new_n470_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT123), .Z(new_n859_));
  NAND2_X1  g658(.A1(new_n834_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n525_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n338_), .ZN(G1344gat));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n582_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n339_), .ZN(G1345gat));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n860_), .B2(new_n631_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n834_), .A2(KEYINPUT124), .A3(new_n680_), .A4(new_n859_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1346gat));
  OAI21_X1  g669(.A(G162gat), .B1(new_n860_), .B2(new_n684_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n611_), .A2(G162gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n860_), .B2(new_n872_), .ZN(G1347gat));
  AOI22_X1  g672(.A1(new_n823_), .A2(new_n631_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n447_), .A2(new_n449_), .A3(new_n490_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n874_), .A2(new_n654_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT126), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n725_), .A3(new_n292_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n874_), .A2(new_n525_), .A3(new_n654_), .A4(new_n876_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n217_), .B1(new_n884_), .B2(KEYINPUT125), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n874_), .A2(new_n654_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n725_), .A3(new_n875_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n885_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n885_), .B2(new_n889_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n883_), .B1(new_n891_), .B2(new_n892_), .ZN(G1348gat));
  NOR3_X1   g692(.A1(new_n878_), .A2(new_n218_), .A3(new_n582_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n882_), .A2(new_n583_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n291_), .ZN(G1349gat));
  AOI21_X1  g695(.A(G183gat), .B1(new_n877_), .B2(new_n680_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n631_), .A2(new_n207_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n882_), .B2(new_n898_), .ZN(G1350gat));
  AND2_X1   g698(.A1(new_n879_), .A2(new_n881_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n636_), .A2(new_n206_), .A3(new_n211_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n684_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n902_));
  OAI22_X1  g701(.A1(new_n900_), .A2(new_n901_), .B1(new_n902_), .B2(new_n204_), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n857_), .A2(new_n449_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n886_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n525_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n237_), .ZN(G1352gat));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n582_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n234_), .ZN(G1353gat));
  AND2_X1   g708(.A1(new_n886_), .A2(new_n904_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n631_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n912_), .B(new_n913_), .Z(G1354gat));
  NAND3_X1  g713(.A1(new_n910_), .A2(new_n245_), .A3(new_n636_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G218gat), .B1(new_n905_), .B2(new_n684_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1355gat));
endmodule


