//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G155gat), .B2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n203_), .B(new_n206_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n203_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n219_));
  XOR2_X1   g018(.A(G155gat), .B(G162gat), .Z(new_n220_));
  AND3_X1   g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n219_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n202_), .B(new_n211_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n220_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT85), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n224_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(new_n202_), .A3(new_n211_), .A4(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G22gat), .B(G50gat), .Z(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT87), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G197gat), .A2(G204gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(KEYINPUT21), .A3(new_n238_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n211_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(KEYINPUT29), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G228gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(G78gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G106gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n248_), .B(new_n252_), .Z(new_n253_));
  OR2_X1    g052(.A1(new_n236_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n235_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT87), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n233_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n236_), .A3(new_n253_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT19), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT24), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR3_X1   g064(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT23), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270_));
  INV_X1    g069(.A(G169gat), .ZN(new_n271_));
  INV_X1    g070(.A(G176gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n273_), .A2(KEYINPUT24), .A3(new_n264_), .A4(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n267_), .A2(new_n269_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT26), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G190gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT88), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(new_n280_), .A3(KEYINPUT88), .ZN(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT25), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G183gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n282_), .A2(new_n283_), .A3(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n268_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n292_), .B2(new_n268_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n274_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT22), .B(G169gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n272_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n276_), .A2(new_n290_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT20), .B1(new_n298_), .B2(new_n246_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT24), .B1(new_n273_), .B2(new_n264_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n268_), .B(new_n292_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT79), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n285_), .A2(new_n287_), .A3(new_n278_), .A4(new_n280_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n275_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n267_), .A2(new_n305_), .A3(new_n269_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT22), .B(G169gat), .Z(new_n308_));
  AND2_X1   g107(.A1(new_n308_), .A2(KEYINPUT80), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n271_), .A2(KEYINPUT22), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n272_), .B1(new_n310_), .B2(KEYINPUT80), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n274_), .B(new_n294_), .C1(new_n309_), .C2(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n246_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n262_), .B1(new_n299_), .B2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G8gat), .B(G36gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n298_), .B2(new_n246_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n307_), .A2(new_n312_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n244_), .A2(new_n245_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n262_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n314_), .A2(new_n319_), .A3(new_n326_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n299_), .A2(new_n313_), .A3(new_n262_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n294_), .A2(new_n297_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n283_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n330_), .A2(new_n281_), .A3(new_n288_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n267_), .A2(new_n269_), .A3(new_n275_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n323_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT94), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT94), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n336_), .B(KEYINPUT20), .C1(new_n333_), .C2(new_n323_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(new_n324_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n328_), .B1(new_n338_), .B2(new_n262_), .ZN(new_n339_));
  OAI211_X1 g138(.A(KEYINPUT27), .B(new_n327_), .C1(new_n339_), .C2(new_n319_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n320_), .B1(new_n333_), .B2(new_n323_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n246_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n325_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT20), .B(new_n325_), .C1(new_n333_), .C2(new_n323_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n246_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n319_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n344_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n319_), .B1(new_n314_), .B2(new_n326_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n341_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n340_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n260_), .A2(new_n353_), .A3(KEYINPUT97), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT97), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n259_), .B2(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G85gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G134gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G127gat), .ZN(new_n367_));
  INV_X1    g166(.A(G127gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G134gat), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n367_), .A2(new_n369_), .A3(KEYINPUT82), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT82), .B1(new_n367_), .B2(new_n369_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n365_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n368_), .A2(G134gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n366_), .A2(G127gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n367_), .A2(new_n369_), .A3(KEYINPUT82), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n364_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n247_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n379_), .B(new_n211_), .C1(new_n222_), .C2(new_n221_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n229_), .A2(KEYINPUT91), .A3(new_n211_), .A4(new_n379_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n363_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n387_), .B(KEYINPUT92), .Z(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n381_), .A2(KEYINPUT4), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n386_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n385_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n362_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(KEYINPUT4), .ZN(new_n396_));
  INV_X1    g195(.A(new_n390_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n388_), .A3(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n361_), .A3(new_n393_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT95), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT81), .B(G43gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n322_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(G15gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT30), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n408_), .A2(new_n412_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT83), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n413_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n379_), .B(KEYINPUT31), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n420_), .ZN(new_n422_));
  OAI211_X1 g221(.A(KEYINPUT83), .B(new_n422_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n357_), .A2(new_n404_), .A3(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n421_), .A2(KEYINPUT84), .A3(new_n423_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT84), .B1(new_n421_), .B2(new_n423_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n399_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n361_), .B1(new_n392_), .B2(new_n388_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n390_), .B1(new_n392_), .B2(KEYINPUT4), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT93), .B1(new_n432_), .B2(new_n389_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  NOR4_X1   g233(.A1(new_n386_), .A2(new_n434_), .A3(new_n388_), .A4(new_n390_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n431_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n398_), .A2(KEYINPUT33), .A3(new_n361_), .A4(new_n393_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT90), .B1(new_n349_), .B2(new_n350_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n348_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n327_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n430_), .A2(new_n436_), .A3(new_n437_), .A4(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n344_), .A2(new_n347_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n339_), .B2(new_n445_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n399_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n361_), .B1(new_n398_), .B2(new_n393_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n259_), .B1(new_n443_), .B2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n340_), .A2(new_n254_), .A3(new_n351_), .A4(new_n258_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n402_), .A2(new_n453_), .A3(new_n403_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n428_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT96), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(new_n428_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n425_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G141gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT77), .ZN(new_n461_));
  XOR2_X1   g260(.A(G169gat), .B(G197gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT76), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G8gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G22gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n410_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G15gat), .A2(G22gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G1gat), .A2(G8gat), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n470_), .A2(new_n471_), .B1(KEYINPUT14), .B2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n468_), .A2(new_n473_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G43gat), .B(G50gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n465_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT75), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n479_), .B(KEYINPUT15), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n476_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n482_), .A3(new_n465_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n464_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n483_), .A2(KEYINPUT75), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n490_));
  AOI211_X1 g289(.A(new_n490_), .B(new_n465_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n464_), .B(new_n487_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n459_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT64), .ZN(new_n496_));
  NAND2_X1  g295(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n496_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT10), .ZN(new_n501_));
  INV_X1    g300(.A(G99gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(KEYINPUT64), .A3(new_n497_), .ZN(new_n504_));
  AOI21_X1  g303(.A(G106gat), .B1(new_n500_), .B2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(KEYINPUT9), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT6), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(G99gat), .A3(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(G85gat), .A3(G92gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n505_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n506_), .A2(new_n507_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n513_), .ZN(new_n521_));
  OR3_X1    g320(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n520_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n523_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n519_), .B1(new_n530_), .B2(new_n513_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n526_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n517_), .A2(new_n527_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT11), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n538_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OR3_X1    g343(.A1(new_n534_), .A2(new_n535_), .A3(new_n544_), .ZN(new_n545_));
  OAI22_X1  g344(.A1(new_n531_), .A2(new_n532_), .B1(new_n505_), .B2(new_n516_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n525_), .A2(new_n526_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n544_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n517_), .A2(new_n527_), .A3(new_n543_), .A4(new_n533_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n535_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n549_), .A2(new_n551_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n544_), .B(new_n555_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n534_), .B2(new_n544_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n554_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G120gat), .B(G148gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n565_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n566_), .A2(KEYINPUT68), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT68), .B1(new_n566_), .B2(new_n567_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n485_), .A2(new_n534_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n575_), .B(new_n578_), .C1(new_n480_), .C2(new_n534_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT69), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n579_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT36), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT37), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n585_), .B(KEYINPUT36), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n582_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n543_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n476_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  XOR2_X1   g395(.A(G127gat), .B(G155gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n595_), .A2(new_n596_), .A3(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT73), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n601_), .B(KEYINPUT17), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT74), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n582_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT70), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n590_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n609_), .B2(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n587_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n592_), .B(new_n607_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n495_), .A2(new_n574_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(G1gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n404_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n612_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n459_), .A2(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n573_), .A2(new_n494_), .A3(new_n607_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n616_), .B1(new_n624_), .B2(new_n617_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n619_), .B2(new_n618_), .ZN(G1324gat));
  INV_X1    g426(.A(G8gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n624_), .B2(new_n352_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT39), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n615_), .A2(new_n628_), .A3(new_n352_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT98), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  INV_X1    g434(.A(new_n428_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n410_), .B1(new_n624_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT41), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n615_), .A2(new_n410_), .A3(new_n636_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1326gat));
  AOI21_X1  g439(.A(new_n469_), .B1(new_n624_), .B2(new_n259_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT42), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n615_), .A2(new_n469_), .A3(new_n259_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1327gat));
  INV_X1    g443(.A(new_n494_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n574_), .A2(new_n645_), .A3(new_n607_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n425_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n403_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(new_n259_), .A3(new_n353_), .A4(new_n401_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n447_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n396_), .A2(new_n389_), .A3(new_n397_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n434_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n432_), .A2(KEYINPUT93), .A3(new_n389_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n654_), .A2(new_n431_), .B1(new_n429_), .B2(new_n399_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n442_), .A2(new_n437_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n650_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n649_), .B1(new_n657_), .B2(new_n259_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n457_), .B1(new_n658_), .B2(new_n428_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n458_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n647_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n592_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n459_), .B2(new_n663_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n646_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n667_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n404_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n607_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n612_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT101), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n495_), .A2(new_n574_), .A3(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n404_), .A2(G29gat), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT102), .Z(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n675_), .A2(new_n682_), .ZN(G1328gat));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n679_), .A2(new_n684_), .A3(new_n352_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT45), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT103), .B(new_n352_), .C1(new_n670_), .C2(new_n673_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G36gat), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n665_), .A2(new_n666_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n646_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n671_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n672_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT103), .B1(new_n696_), .B2(new_n352_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n686_), .B1(new_n688_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT46), .B(new_n686_), .C1(new_n688_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n679_), .A2(new_n703_), .A3(new_n636_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n424_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n674_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n706_), .B2(new_n703_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT47), .B(new_n704_), .C1(new_n706_), .C2(new_n703_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n679_), .B2(new_n259_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n259_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n696_), .B2(new_n713_), .ZN(G1331gat));
  NAND4_X1  g513(.A1(new_n622_), .A2(new_n494_), .A3(new_n573_), .A4(new_n676_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n404_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n573_), .A2(new_n494_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n459_), .A2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n614_), .ZN(new_n719_));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n617_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n715_), .B2(new_n353_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n719_), .A2(new_n725_), .A3(new_n352_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n715_), .B2(new_n428_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n719_), .A2(new_n730_), .A3(new_n636_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1334gat));
  OAI21_X1  g531(.A(G78gat), .B1(new_n715_), .B2(new_n260_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT50), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n719_), .A2(new_n250_), .A3(new_n259_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1335gat));
  INV_X1    g535(.A(new_n689_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT105), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(KEYINPUT105), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n717_), .A2(new_n676_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n404_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n718_), .A2(new_n678_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT104), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT104), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(G85gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n617_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n742_), .A2(new_n748_), .ZN(G1336gat));
  AOI21_X1  g548(.A(G92gat), .B1(new_n746_), .B2(new_n352_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT106), .ZN(new_n751_));
  INV_X1    g550(.A(G92gat), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n741_), .A2(new_n752_), .A3(new_n353_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n741_), .B2(new_n428_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n705_), .B1(new_n504_), .B2(new_n500_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT51), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(new_n759_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1338gat));
  NAND2_X1  g563(.A1(new_n740_), .A2(new_n259_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G106gat), .B1(new_n737_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT52), .ZN(new_n767_));
  INV_X1    g566(.A(G106gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n746_), .A2(new_n768_), .A3(new_n259_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g570(.A(new_n465_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n486_), .A2(new_n482_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n463_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n484_), .A2(new_n487_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n463_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n567_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n548_), .A2(KEYINPUT12), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n556_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n549_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n552_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n559_), .A2(KEYINPUT55), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n780_), .B2(new_n554_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n565_), .ZN(new_n789_));
  OAI211_X1 g588(.A(KEYINPUT108), .B(new_n782_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n789_), .A4(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n559_), .A2(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n780_), .A2(new_n784_), .A3(new_n554_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n792_), .A2(new_n793_), .B1(new_n552_), .B2(new_n781_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n565_), .B1(new_n794_), .B2(KEYINPUT108), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n788_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n796_), .B2(KEYINPUT110), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n789_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n792_), .A2(new_n793_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT108), .B1(new_n800_), .B2(new_n782_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n798_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT58), .B(new_n778_), .C1(new_n797_), .C2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n778_), .B1(new_n797_), .B2(new_n804_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n663_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n777_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n567_), .B1(new_n488_), .B2(new_n493_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n802_), .B2(new_n791_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(KEYINPUT109), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n813_), .B(new_n810_), .C1(new_n802_), .C2(new_n791_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n612_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n805_), .A2(new_n808_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT57), .B(new_n612_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n676_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n574_), .A2(new_n614_), .A3(new_n494_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n819_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n357_), .A2(new_n617_), .A3(new_n424_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n645_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n815_), .A2(new_n816_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n806_), .A2(new_n807_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n664_), .A3(new_n805_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(new_n832_), .A3(KEYINPUT112), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n818_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n822_), .B1(new_n837_), .B2(new_n607_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT111), .B(KEYINPUT59), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n824_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT113), .B1(new_n829_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843_));
  OAI221_X1 g642(.A(new_n843_), .B1(new_n838_), .B2(new_n840_), .C1(new_n828_), .C2(new_n825_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n842_), .A2(new_n844_), .A3(new_n645_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n827_), .B1(new_n845_), .B2(new_n826_), .ZN(G1340gat));
  XOR2_X1   g645(.A(KEYINPUT114), .B(G120gat), .Z(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n574_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n825_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT115), .Z(new_n850_));
  OR3_X1    g649(.A1(new_n829_), .A2(new_n841_), .A3(new_n574_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n847_), .B2(new_n852_), .ZN(G1341gat));
  NAND3_X1  g652(.A1(new_n825_), .A2(new_n368_), .A3(new_n676_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n842_), .A2(new_n844_), .A3(new_n676_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n368_), .ZN(G1342gat));
  NAND3_X1  g655(.A1(new_n825_), .A2(new_n366_), .A3(new_n621_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n842_), .A2(new_n844_), .A3(new_n664_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n366_), .ZN(G1343gat));
  NOR3_X1   g658(.A1(new_n636_), .A2(new_n404_), .A3(new_n453_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT116), .B1(new_n823_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n860_), .C1(new_n819_), .C2(new_n822_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n645_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n573_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT117), .B(G148gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n676_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT118), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n865_), .A2(new_n873_), .A3(new_n676_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n872_), .A2(new_n874_), .A3(new_n876_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n865_), .A2(new_n881_), .A3(new_n621_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n663_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT119), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n882_), .B(new_n886_), .C1(new_n881_), .C2(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1347gat));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n617_), .A2(new_n353_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n636_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n259_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n645_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT120), .B1(new_n838_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895_));
  INV_X1    g694(.A(new_n893_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n818_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n676_), .B1(new_n898_), .B2(new_n836_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n895_), .B(new_n896_), .C1(new_n899_), .C2(new_n822_), .ZN(new_n900_));
  AND2_X1   g699(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n894_), .A2(G169gat), .A3(new_n900_), .A4(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n892_), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT122), .B1(new_n838_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n892_), .C1(new_n899_), .C2(new_n822_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n494_), .A2(new_n308_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n902_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n901_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n818_), .B1(new_n817_), .B2(KEYINPUT112), .ZN(new_n913_));
  INV_X1    g712(.A(new_n836_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n607_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n822_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n893_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n271_), .B1(new_n917_), .B2(new_n895_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n912_), .B1(new_n918_), .B2(new_n894_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n889_), .B1(new_n909_), .B2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n894_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n900_), .A2(G169gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n911_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n923_), .A2(KEYINPUT123), .A3(new_n902_), .A4(new_n908_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n924_), .ZN(G1348gat));
  NAND3_X1  g724(.A1(new_n904_), .A2(new_n573_), .A3(new_n906_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n272_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT124), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n926_), .A2(new_n929_), .A3(new_n272_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n823_), .A2(new_n259_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n574_), .A2(new_n891_), .A3(new_n272_), .ZN(new_n932_));
  AOI22_X1  g731(.A1(new_n928_), .A2(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  AND2_X1   g732(.A1(new_n904_), .A2(new_n906_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n607_), .A2(new_n289_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n931_), .A2(new_n636_), .A3(new_n676_), .A4(new_n890_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n934_), .A2(new_n935_), .B1(new_n284_), .B2(new_n936_), .ZN(G1350gat));
  NAND4_X1  g736(.A1(new_n934_), .A2(new_n282_), .A3(new_n283_), .A4(new_n621_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n904_), .A2(new_n664_), .A3(new_n906_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n939_), .A2(new_n940_), .A3(G190gat), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n939_), .B2(G190gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n938_), .B1(new_n941_), .B2(new_n942_), .ZN(G1351gat));
  NAND3_X1  g742(.A1(new_n890_), .A2(new_n259_), .A3(new_n428_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n823_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n645_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT126), .B(G197gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n946_), .B(new_n947_), .ZN(G1352gat));
  NAND2_X1  g747(.A1(new_n945_), .A2(new_n573_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n949_), .B(new_n950_), .Z(G1353gat));
  NAND2_X1  g750(.A1(new_n945_), .A2(new_n676_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  AND2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n952_), .A2(new_n953_), .A3(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n952_), .B2(new_n953_), .ZN(G1354gat));
  INV_X1    g755(.A(G218gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n945_), .A2(new_n957_), .A3(new_n621_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n823_), .A2(new_n663_), .A3(new_n944_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n957_), .ZN(G1355gat));
endmodule


