//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT80), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT31), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n202_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(new_n207_), .B2(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G227gat), .A2(G233gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT78), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT30), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT23), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n216_), .A2(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT25), .B(G183gat), .ZN(new_n226_));
  INV_X1    g025(.A(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT26), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT26), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n227_), .A2(KEYINPUT77), .A3(KEYINPUT26), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n226_), .A2(new_n230_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n225_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G169gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n215_), .A2(new_n217_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n238_), .B(new_n239_), .C1(G183gat), .C2(G190gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G71gat), .B(G99gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(G15gat), .B(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n242_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n209_), .A2(new_n213_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n214_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n246_), .B1(new_n214_), .B2(new_n247_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n256_), .A2(new_n259_), .A3(new_n252_), .A4(new_n257_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G197gat), .B(G204gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n251_), .B1(new_n265_), .B2(new_n252_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT88), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G218gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(G211gat), .ZN(new_n269_));
  INV_X1    g068(.A(G211gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G218gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n258_), .A2(G197gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n257_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(KEYINPUT21), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n263_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n262_), .B1(new_n267_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT86), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(G228gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(G228gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287_));
  INV_X1    g086(.A(G155gat), .ZN(new_n288_));
  INV_X1    g087(.A(G162gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT1), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G155gat), .A3(G162gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n290_), .A2(new_n292_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G141gat), .ZN(new_n297_));
  INV_X1    g096(.A(G148gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n286_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n296_), .A2(new_n286_), .A3(new_n301_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n290_), .A2(new_n295_), .A3(new_n291_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT84), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT84), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n290_), .A2(new_n308_), .A3(new_n295_), .A4(new_n291_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n299_), .A2(KEYINPUT3), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n299_), .A2(KEYINPUT3), .B1(new_n312_), .B2(new_n300_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n314_), .A2(KEYINPUT83), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(KEYINPUT83), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n311_), .B(new_n313_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n310_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n310_), .A2(new_n317_), .A3(KEYINPUT85), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n305_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n285_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n304_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(new_n302_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n310_), .A2(KEYINPUT85), .A3(new_n317_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT85), .B1(new_n310_), .B2(new_n317_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n330_));
  AOI21_X1  g129(.A(new_n278_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n284_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n324_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G78gat), .B(G106gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n324_), .B(new_n336_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT90), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n322_), .A2(new_n323_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT28), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n341_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n338_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n335_), .A2(new_n344_), .A3(new_n339_), .A4(new_n337_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n205_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT94), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n322_), .B2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n350_), .B(new_n326_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(new_n205_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT4), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OR3_X1    g155(.A1(new_n322_), .A2(KEYINPUT4), .A3(new_n205_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n352_), .B(new_n205_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n355_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT95), .B(G85gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT0), .B(G57gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n358_), .A2(KEYINPUT33), .A3(new_n360_), .A4(new_n366_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n276_), .B1(new_n275_), .B2(new_n263_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n255_), .A2(G204gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n258_), .A2(G197gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT21), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  AND4_X1   g173(.A1(new_n276_), .A2(new_n263_), .A3(new_n374_), .A4(new_n251_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n261_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT26), .B(G190gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n226_), .A2(new_n377_), .B1(new_n379_), .B2(new_n223_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n221_), .B1(new_n380_), .B2(KEYINPUT91), .ZN(new_n381_));
  XOR2_X1   g180(.A(KEYINPUT25), .B(G183gat), .Z(new_n382_));
  NAND2_X1  g181(.A1(new_n232_), .A2(new_n228_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n224_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT91), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n241_), .B1(new_n381_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT92), .B1(new_n376_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n376_), .B2(new_n242_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n241_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n221_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n380_), .A2(KEYINPUT91), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n278_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n388_), .A2(new_n390_), .A3(new_n393_), .A4(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n398_), .B2(new_n278_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n376_), .A2(new_n242_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n392_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n407_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n401_), .A2(new_n404_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT93), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n401_), .A2(new_n404_), .A3(new_n414_), .A4(new_n411_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n401_), .A2(new_n404_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n410_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n413_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n366_), .B1(new_n359_), .B2(new_n356_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n369_), .A2(new_n370_), .A3(new_n418_), .A4(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n408_), .A2(KEYINPUT32), .A3(new_n409_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n389_), .B1(new_n376_), .B2(new_n387_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n425_), .B(new_n393_), .C1(new_n376_), .C2(new_n242_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n394_), .B1(new_n234_), .B2(new_n225_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n278_), .B2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n376_), .A2(new_n387_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n392_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n424_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n423_), .B(KEYINPUT96), .ZN(new_n433_));
  OAI22_X1  g232(.A1(new_n431_), .A2(new_n432_), .B1(new_n416_), .B2(new_n433_), .ZN(new_n434_));
  AOI211_X1 g233(.A(KEYINPUT97), .B(new_n424_), .C1(new_n426_), .C2(new_n430_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n358_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n366_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n348_), .B1(new_n422_), .B2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n437_), .A2(new_n438_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n413_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n426_), .A2(new_n430_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n410_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n412_), .A2(KEYINPUT27), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n442_), .A2(new_n443_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n441_), .A2(new_n348_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n250_), .B1(new_n440_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT98), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT98), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n250_), .C1(new_n440_), .C2(new_n448_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n441_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(new_n250_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n442_), .A2(new_n443_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n446_), .A2(new_n445_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n457_), .A2(new_n348_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n330_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n376_), .B1(new_n322_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n461_), .A2(new_n284_), .B1(new_n462_), .B2(new_n285_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT90), .B1(new_n463_), .B2(new_n336_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n464_), .A2(new_n344_), .B1(new_n337_), .B2(new_n335_), .ZN(new_n465_));
  AND4_X1   g264(.A1(new_n339_), .A2(new_n335_), .A3(new_n337_), .A4(new_n344_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT99), .B1(new_n467_), .B2(new_n447_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n454_), .B1(new_n459_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT100), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT100), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n454_), .B(new_n471_), .C1(new_n459_), .C2(new_n468_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n450_), .A2(new_n452_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n477_), .B1(KEYINPUT65), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(new_n477_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n476_), .B1(new_n481_), .B2(KEYINPUT66), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(KEYINPUT66), .B2(new_n481_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G85gat), .B(G92gat), .Z(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(KEYINPUT8), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n481_), .B2(new_n476_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT8), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT10), .B(G99gat), .Z(new_n490_));
  AOI21_X1  g289(.A(new_n476_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(KEYINPUT64), .ZN(new_n492_));
  INV_X1    g291(.A(G85gat), .ZN(new_n493_));
  INV_X1    g292(.A(G92gat), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT9), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n484_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n488_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n485_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G29gat), .B(G36gat), .Z(new_n501_));
  XOR2_X1   g300(.A(G43gat), .B(G50gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n500_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n485_), .A2(new_n499_), .A3(new_n507_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(KEYINPUT35), .A3(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n510_), .A2(new_n518_), .A3(new_n511_), .A4(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G190gat), .B(G218gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G134gat), .B(G162gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n523_), .B(KEYINPUT36), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n523_), .A2(KEYINPUT36), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n517_), .A2(new_n526_), .A3(new_n519_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n473_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G71gat), .B(G78gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT11), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(new_n535_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n500_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n485_), .A2(new_n499_), .A3(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(KEYINPUT67), .A3(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(KEYINPUT12), .A3(new_n543_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n500_), .A2(new_n553_), .A3(new_n541_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n546_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n533_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n545_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n533_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n558_), .A2(new_n549_), .A3(new_n550_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT13), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT13), .B1(new_n556_), .B2(new_n560_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT76), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G15gat), .B(G22gat), .ZN(new_n567_));
  INV_X1    g366(.A(G1gat), .ZN(new_n568_));
  INV_X1    g367(.A(G8gat), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT14), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G1gat), .B(G8gat), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n572_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n507_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT72), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n509_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT73), .ZN(new_n581_));
  INV_X1    g380(.A(new_n507_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n577_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT73), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n575_), .A2(KEYINPUT72), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n575_), .A2(KEYINPUT72), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n588_), .A2(new_n589_), .B1(new_n509_), .B2(new_n578_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n587_), .B1(new_n590_), .B2(new_n577_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n581_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G113gat), .B(G141gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT74), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT75), .B(new_n566_), .C1(new_n592_), .C2(new_n596_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n588_), .A2(new_n589_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n580_), .B(KEYINPUT73), .C1(new_n577_), .C2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n590_), .A2(new_n587_), .A3(new_n577_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT76), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n600_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n596_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n597_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n597_), .B2(new_n603_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n565_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n578_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n541_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(KEYINPUT71), .A2(KEYINPUT17), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n614_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  MUX2_X1   g419(.A(new_n619_), .B(KEYINPUT17), .S(new_n618_), .Z(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n610_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n529_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n453_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n568_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  INV_X1    g428(.A(new_n609_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n473_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n525_), .A2(KEYINPUT70), .A3(new_n527_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n525_), .A2(KEYINPUT70), .A3(KEYINPUT37), .A4(new_n527_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n623_), .A3(new_n635_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n631_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n568_), .A3(new_n453_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n628_), .B1(new_n629_), .B2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n629_), .B2(new_n640_), .ZN(G1324gat));
  NAND3_X1  g441(.A1(new_n529_), .A2(new_n457_), .A3(new_n625_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT101), .A3(G8gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT101), .B1(new_n643_), .B2(G8gat), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n447_), .A2(G8gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g452(.A(G15gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n250_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n626_), .B2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT41), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n639_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n626_), .B2(new_n348_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT42), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n639_), .A2(new_n660_), .A3(new_n348_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n610_), .A2(new_n623_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n450_), .A2(new_n452_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n470_), .A2(new_n472_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n634_), .A2(new_n635_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n673_));
  INV_X1    g472(.A(new_n671_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n473_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n666_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n669_), .A2(new_n671_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT103), .B1(new_n677_), .B2(new_n673_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT44), .B(new_n665_), .C1(new_n676_), .C2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n453_), .A2(G29gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n665_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n673_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT43), .B(new_n674_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT103), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n675_), .A2(new_n666_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n681_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n679_), .B(new_n680_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n565_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n528_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n623_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n631_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G29gat), .B1(new_n696_), .B2(new_n453_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n690_), .A2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT105), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT106), .Z(new_n701_));
  OAI211_X1 g500(.A(new_n457_), .B(new_n679_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G36gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n699_), .A2(KEYINPUT105), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n447_), .A2(G36gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n696_), .B2(new_n706_), .ZN(new_n707_));
  AND4_X1   g506(.A1(new_n705_), .A2(new_n631_), .A3(new_n695_), .A4(new_n706_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n701_), .B1(new_n703_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n701_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n712_), .B(new_n709_), .C1(new_n702_), .C2(G36gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1329gat));
  INV_X1    g513(.A(G43gat), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n250_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n679_), .B(new_n716_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n696_), .A2(new_n655_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT47), .ZN(G1330gat));
  AND2_X1   g520(.A1(new_n348_), .A2(G50gat), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n679_), .B(new_n722_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G50gat), .B1(new_n696_), .B2(new_n348_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n691_), .A2(new_n630_), .ZN(new_n727_));
  NOR4_X1   g526(.A1(new_n473_), .A2(new_n624_), .A3(new_n528_), .A4(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(G57gat), .A3(new_n453_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n729_), .A2(new_n730_), .ZN(new_n732_));
  NOR4_X1   g531(.A1(new_n473_), .A2(new_n609_), .A3(new_n565_), .A4(new_n636_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n453_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(G1332gat));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n728_), .B2(new_n457_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT48), .Z(new_n738_));
  NAND2_X1  g537(.A1(new_n457_), .A2(new_n736_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT108), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n733_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n728_), .B2(new_n655_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT49), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n733_), .A2(new_n743_), .A3(new_n655_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  INV_X1    g546(.A(G78gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n728_), .B2(new_n348_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT50), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n748_), .A3(new_n348_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1335gat));
  NOR4_X1   g551(.A1(new_n473_), .A2(new_n609_), .A3(new_n565_), .A4(new_n694_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT109), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n493_), .A3(new_n453_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n685_), .A2(new_n686_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n727_), .A2(new_n623_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n453_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n759_), .B2(new_n493_), .ZN(G1336gat));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n494_), .A3(new_n457_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n457_), .A3(new_n757_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n763_), .B2(new_n494_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n655_), .A3(new_n490_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n655_), .B(new_n757_), .C1(new_n676_), .C2(new_n678_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G99gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G99gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n765_), .B(new_n772_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n754_), .A2(new_n489_), .A3(new_n348_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n348_), .B(new_n757_), .C1(new_n676_), .C2(new_n678_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G106gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n775_), .B(new_n782_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  NOR2_X1   g583(.A1(new_n459_), .A2(new_n468_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n655_), .A2(new_n453_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n791_));
  INV_X1    g590(.A(new_n560_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n607_), .A2(new_n608_), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n552_), .A2(new_n546_), .A3(new_n554_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n558_), .A2(KEYINPUT55), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n559_), .B1(new_n555_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT112), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(KEYINPUT111), .A3(new_n799_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT112), .B1(new_n799_), .B2(KEYINPUT111), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n795_), .A2(new_n797_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n590_), .A2(new_n585_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n596_), .C1(new_n585_), .C2(new_n598_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT113), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n584_), .A2(new_n577_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n805_), .A3(new_n809_), .A4(new_n596_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n601_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n793_), .A2(new_n804_), .B1(new_n561_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n791_), .B1(new_n813_), .B2(new_n528_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n798_), .B(new_n799_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n792_), .A2(new_n601_), .A3(new_n811_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n798_), .A2(new_n799_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n797_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n816_), .B(KEYINPUT58), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n671_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n814_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n561_), .A2(new_n812_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n800_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n608_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n597_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n560_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n692_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n824_), .A2(KEYINPUT117), .B1(new_n832_), .B2(KEYINPUT57), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n814_), .A2(new_n834_), .A3(new_n823_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n623_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n637_), .B2(new_n630_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n636_), .ZN(new_n839_));
  AND4_X1   g638(.A1(new_n837_), .A2(new_n565_), .A3(new_n630_), .A4(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n790_), .B1(new_n836_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n822_), .A2(new_n671_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT58), .B1(new_n815_), .B2(new_n816_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n831_), .B2(new_n791_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n830_), .A2(KEYINPUT57), .A3(new_n692_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n623_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n787_), .B1(new_n849_), .B2(new_n841_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n843_), .B1(new_n850_), .B2(KEYINPUT59), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n814_), .A2(new_n848_), .A3(new_n823_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n841_), .B1(new_n852_), .B2(new_n624_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n843_), .B(KEYINPUT59), .C1(new_n853_), .C2(new_n788_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n842_), .B1(new_n851_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n630_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n630_), .A2(G113gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n850_), .B2(new_n858_), .ZN(G1340gat));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n856_), .B2(new_n565_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT59), .B1(new_n853_), .B2(new_n788_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT115), .ZN(new_n863_));
  INV_X1    g662(.A(new_n791_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n830_), .B2(new_n692_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT117), .B1(new_n865_), .B2(new_n846_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n848_), .A3(new_n835_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n624_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n841_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n863_), .A2(new_n854_), .B1(new_n870_), .B2(new_n790_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(KEYINPUT118), .A3(new_n691_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n861_), .A2(G120gat), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n850_), .ZN(new_n874_));
  INV_X1    g673(.A(G120gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n565_), .B2(KEYINPUT60), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n874_), .B(new_n876_), .C1(KEYINPUT60), .C2(new_n875_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(G1341gat));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879_));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n871_), .B2(new_n623_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n850_), .A2(G127gat), .A3(new_n624_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n623_), .B(new_n842_), .C1(new_n851_), .C2(new_n855_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G127gat), .ZN(new_n885_));
  INV_X1    g684(.A(new_n882_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(KEYINPUT119), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(G1342gat));
  OAI21_X1  g687(.A(G134gat), .B1(new_n856_), .B2(new_n674_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n692_), .A2(G134gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n850_), .B2(new_n890_), .ZN(G1343gat));
  NOR4_X1   g690(.A1(new_n655_), .A2(new_n467_), .A3(new_n457_), .A4(new_n441_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n853_), .A2(KEYINPUT120), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT120), .B1(new_n853_), .B2(new_n893_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n609_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n691_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT121), .B(G148gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1345gat));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n897_), .B2(new_n623_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI211_X1 g704(.A(KEYINPUT122), .B(new_n624_), .C1(new_n895_), .C2(new_n896_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT61), .B(G155gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n905_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n908_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1346gat));
  NAND2_X1  g711(.A1(new_n671_), .A2(G162gat), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT123), .Z(new_n914_));
  NAND2_X1  g713(.A1(new_n897_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n692_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(G162gat), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n915_), .B(KEYINPUT124), .C1(G162gat), .C2(new_n916_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n454_), .A2(new_n457_), .ZN(new_n922_));
  AOI211_X1 g721(.A(new_n348_), .B(new_n922_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n609_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n924_), .A2(new_n925_), .A3(G169gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(G169gat), .ZN(new_n927_));
  INV_X1    g726(.A(new_n923_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT22), .B(G169gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n609_), .A2(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT125), .ZN(new_n931_));
  OAI22_X1  g730(.A1(new_n926_), .A2(new_n927_), .B1(new_n928_), .B2(new_n931_), .ZN(G1348gat));
  AOI21_X1  g731(.A(G176gat), .B1(new_n923_), .B2(new_n691_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n853_), .A2(new_n348_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n922_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n691_), .A2(new_n935_), .A3(G176gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n934_), .B2(new_n936_), .ZN(G1349gat));
  NOR2_X1   g736(.A1(new_n624_), .A2(new_n226_), .ZN(new_n938_));
  INV_X1    g737(.A(G183gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n934_), .A2(new_n623_), .A3(new_n935_), .ZN(new_n940_));
  AOI22_X1  g739(.A1(new_n923_), .A2(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n928_), .B2(new_n674_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n923_), .A2(new_n377_), .A3(new_n528_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1351gat));
  INV_X1    g743(.A(new_n853_), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n655_), .A2(new_n453_), .A3(new_n467_), .A4(new_n447_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  AOI22_X1  g747(.A1(new_n948_), .A2(new_n609_), .B1(KEYINPUT126), .B2(G197gat), .ZN(new_n949_));
  NOR2_X1   g748(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n950_), .B(KEYINPUT127), .Z(new_n951_));
  XNOR2_X1  g750(.A(new_n949_), .B(new_n951_), .ZN(G1352gat));
  NOR2_X1   g751(.A1(new_n947_), .A2(new_n565_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(new_n258_), .ZN(G1353gat));
  NAND2_X1  g753(.A1(new_n948_), .A2(new_n623_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  AND2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(new_n955_), .B2(new_n956_), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n947_), .B2(new_n674_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n528_), .A2(new_n268_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n947_), .B2(new_n961_), .ZN(G1355gat));
endmodule


