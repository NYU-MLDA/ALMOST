//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT91), .Z(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT89), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(new_n207_), .B2(new_n204_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT90), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT3), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n203_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n206_), .A2(new_n214_), .ZN(new_n215_));
  OAI221_X1 g014(.A(new_n215_), .B1(KEYINPUT1), .B2(new_n202_), .C1(G141gat), .C2(G148gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G113gat), .B(G120gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n219_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT88), .B1(new_n218_), .B2(new_n219_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n220_), .B(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n224_), .B2(new_n217_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT4), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n213_), .A2(new_n216_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n224_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT101), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n230_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n225_), .A2(new_n234_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G57gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n238_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT102), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G183gat), .ZN(new_n250_));
  INV_X1    g049(.A(G190gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT23), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT83), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(G183gat), .A3(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT84), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(G183gat), .B2(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT22), .B(G169gat), .Z(new_n260_));
  OAI211_X1 g059(.A(new_n258_), .B(new_n259_), .C1(G176gat), .C2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT82), .Z(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n252_), .A2(new_n255_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n266_), .A2(new_n267_), .B1(new_n268_), .B2(new_n262_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n261_), .A2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G211gat), .B(G218gat), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT95), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT21), .ZN(new_n275_));
  AOI211_X1 g074(.A(new_n274_), .B(new_n275_), .C1(G197gat), .C2(G204gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT94), .ZN(new_n277_));
  INV_X1    g076(.A(G197gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n273_), .B(new_n276_), .C1(G204gat), .C2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G204gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G197gat), .ZN(new_n282_));
  OAI221_X1 g081(.A(new_n282_), .B1(new_n281_), .B2(new_n279_), .C1(new_n272_), .C2(new_n275_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n278_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n280_), .A2(new_n283_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n271_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT97), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT26), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT81), .B1(new_n291_), .B2(G190gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT80), .B(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n294_), .A2(KEYINPUT25), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n296_));
  OAI221_X1 g095(.A(new_n292_), .B1(KEYINPUT81), .B2(new_n266_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n263_), .A2(KEYINPUT24), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n297_), .A2(new_n257_), .A3(new_n298_), .A4(new_n264_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n265_), .B1(new_n294_), .B2(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(G176gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(KEYINPUT85), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G169gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(G169gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n286_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n290_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n289_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n287_), .A2(new_n288_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n249_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n271_), .A2(new_n286_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n307_), .B2(new_n308_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n249_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT99), .B(G8gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G36gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n319_), .B(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT100), .B1(new_n316_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n312_), .A2(new_n315_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(KEYINPUT100), .A3(new_n325_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n225_), .A2(new_n234_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n243_), .B(new_n330_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n243_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT33), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n325_), .A2(KEYINPUT32), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n324_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n249_), .B1(new_n287_), .B2(new_n309_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n313_), .A2(new_n314_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n249_), .B2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n244_), .B(new_n337_), .C1(new_n340_), .C2(new_n336_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n224_), .B(KEYINPUT30), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n307_), .B(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G71gat), .B(G99gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT31), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n344_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G15gat), .B(G43gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n352_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT28), .ZN(new_n358_));
  XOR2_X1   g157(.A(G22gat), .B(G50gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n286_), .B1(new_n227_), .B2(KEYINPUT29), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT93), .B(G233gat), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(G228gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n361_), .B(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n366_), .A2(KEYINPUT92), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n360_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n360_), .A2(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n342_), .A2(new_n356_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n327_), .A2(new_n373_), .A3(new_n328_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n326_), .B(KEYINPUT27), .C1(new_n325_), .C2(new_n340_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n356_), .A2(new_n370_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(new_n355_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n245_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n372_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G134gat), .B(G162gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G218gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT73), .B(G190gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT36), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G232gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT34), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT35), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT72), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G85gat), .B(G92gat), .Z(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n397_));
  INV_X1    g196(.A(G99gat), .ZN(new_n398_));
  INV_X1    g197(.A(G106gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT7), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G99gat), .A2(G106gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(KEYINPUT68), .A3(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n407_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n396_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT8), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT69), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n406_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT66), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n407_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT66), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n403_), .A2(new_n423_), .A3(new_n424_), .A4(new_n410_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n420_), .A2(new_n416_), .A3(new_n395_), .A4(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT67), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n412_), .A2(new_n413_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(new_n408_), .A3(new_n403_), .A4(new_n410_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n395_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT8), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n403_), .A2(new_n423_), .A3(new_n410_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT8), .B1(new_n434_), .B2(KEYINPUT66), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n435_), .A2(KEYINPUT67), .A3(new_n395_), .A4(new_n425_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n417_), .A2(new_n428_), .A3(new_n433_), .A4(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G29gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G43gat), .B(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT64), .B1(new_n396_), .B2(KEYINPUT9), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n240_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(KEYINPUT9), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT10), .B(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n412_), .B1(new_n446_), .B2(new_n399_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n437_), .A2(new_n440_), .A3(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n391_), .A2(KEYINPUT35), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n440_), .B(KEYINPUT15), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n437_), .B2(new_n449_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n394_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n455_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n457_), .A2(new_n393_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n389_), .B1(new_n459_), .B2(KEYINPUT74), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(KEYINPUT74), .A3(new_n389_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT75), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465_));
  INV_X1    g264(.A(new_n459_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n386_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(KEYINPUT36), .A3(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470_));
  AOI211_X1 g269(.A(new_n470_), .B(new_n388_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n468_), .B1(new_n460_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT75), .A2(KEYINPUT37), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n465_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n382_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G176gat), .B(G204gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G120gat), .B(G148gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n483_), .A2(KEYINPUT11), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(KEYINPUT11), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G71gat), .B(G78gat), .ZN(new_n486_));
  OR3_X1    g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n486_), .A3(KEYINPUT11), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n437_), .B2(new_n449_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT70), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G230gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n437_), .A2(new_n449_), .A3(new_n489_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n491_), .B(new_n493_), .C1(new_n496_), .C2(new_n490_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n437_), .A2(new_n449_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n489_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT12), .A3(new_n494_), .ZN(new_n502_));
  AOI211_X1 g301(.A(KEYINPUT12), .B(new_n489_), .C1(new_n437_), .C2(new_n449_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n493_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n482_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(KEYINPUT12), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n490_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n492_), .B1(new_n508_), .B2(new_n503_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n482_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n497_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n506_), .A2(KEYINPUT13), .A3(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n489_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G15gat), .B(G22gat), .Z(new_n519_));
  NAND2_X1  g318(.A1(G1gat), .A2(G8gat), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(KEYINPUT14), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT76), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n520_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G1gat), .A2(G8gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n521_), .B(KEYINPUT76), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n518_), .B(new_n531_), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G183gat), .B(G211gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G127gat), .B(G155gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  OR3_X1    g338(.A1(new_n533_), .A2(new_n534_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(KEYINPUT17), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n533_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n516_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n523_), .A2(new_n527_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n529_), .A2(new_n526_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n453_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n528_), .A2(new_n530_), .A3(new_n440_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT78), .ZN(new_n551_));
  INV_X1    g350(.A(new_n548_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n549_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n440_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT78), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n547_), .A2(new_n556_), .A3(new_n549_), .A4(new_n548_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT79), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n560_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n544_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n246_), .B1(new_n477_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n382_), .A2(KEYINPUT102), .A3(new_n568_), .A4(new_n476_), .ZN(new_n569_));
  AOI211_X1 g368(.A(G1gat), .B(new_n245_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT104), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n570_), .A2(new_n571_), .A3(KEYINPUT38), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(KEYINPUT38), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n570_), .B2(KEYINPUT38), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n472_), .B(KEYINPUT103), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n372_), .B2(new_n381_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n577_), .A2(new_n568_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n579_), .B2(new_n245_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .A4(new_n580_), .ZN(G1324gat));
  INV_X1    g380(.A(KEYINPUT40), .ZN(new_n582_));
  AOI21_X1  g381(.A(G8gat), .B1(new_n567_), .B2(new_n569_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n376_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT105), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(KEYINPUT106), .A3(new_n376_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n577_), .A2(new_n568_), .A3(new_n376_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT106), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(G8gat), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n582_), .B1(new_n585_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT105), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n584_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n590_), .B(KEYINPUT39), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(KEYINPUT40), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(G1325gat));
  INV_X1    g397(.A(G15gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n578_), .B2(new_n355_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT41), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n477_), .A2(new_n566_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n599_), .A3(new_n355_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(G1326gat));
  INV_X1    g403(.A(G22gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n578_), .B2(new_n370_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT42), .Z(new_n607_));
  NAND3_X1  g406(.A1(new_n602_), .A2(new_n605_), .A3(new_n370_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1327gat));
  INV_X1    g408(.A(KEYINPUT43), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n469_), .A2(new_n475_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n382_), .B2(new_n611_), .ZN(new_n612_));
  AOI211_X1 g411(.A(KEYINPUT43), .B(new_n476_), .C1(new_n372_), .C2(new_n381_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n560_), .B(new_n563_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n516_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n614_), .A2(KEYINPUT44), .A3(new_n543_), .A4(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n543_), .B(new_n616_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n620_), .A3(new_n244_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT107), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT107), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(G29gat), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n472_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n372_), .B2(new_n381_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n543_), .A3(new_n616_), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n627_), .A2(G29gat), .A3(new_n245_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(G1328gat));
  NAND3_X1  g428(.A1(new_n617_), .A2(new_n620_), .A3(new_n376_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G36gat), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT45), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n627_), .A2(G36gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n376_), .B(KEYINPUT108), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  OR4_X1    g434(.A1(new_n632_), .A2(new_n627_), .A3(G36gat), .A4(new_n634_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n631_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT46), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n631_), .A2(new_n637_), .A3(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1329gat));
  NAND3_X1  g441(.A1(new_n617_), .A2(new_n620_), .A3(new_n355_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G43gat), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n627_), .A2(G43gat), .A3(new_n356_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT47), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(KEYINPUT47), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1330gat));
  NAND3_X1  g449(.A1(new_n617_), .A2(new_n620_), .A3(new_n370_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G50gat), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n371_), .A2(G50gat), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT109), .Z(new_n654_));
  OR2_X1    g453(.A1(new_n627_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT110), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(KEYINPUT110), .A3(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1331gat));
  INV_X1    g459(.A(new_n516_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n565_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n477_), .A2(new_n543_), .A3(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT111), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT111), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n244_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G57gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n663_), .A2(new_n543_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n577_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n245_), .A2(new_n668_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n667_), .A2(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(G1332gat));
  INV_X1    g471(.A(G64gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n634_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n664_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n670_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G64gat), .B1(new_n676_), .B2(new_n634_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT48), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT48), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT112), .ZN(G1333gat));
  INV_X1    g480(.A(G71gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n670_), .B2(new_n355_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n664_), .A2(new_n682_), .A3(new_n355_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1334gat));
  INV_X1    g486(.A(G78gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n670_), .B2(new_n370_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT50), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n664_), .A2(new_n688_), .A3(new_n370_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1335gat));
  NAND3_X1  g491(.A1(new_n626_), .A2(new_n543_), .A3(new_n662_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n614_), .A2(new_n543_), .A3(new_n662_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT114), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(KEYINPUT114), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n245_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n699_), .B2(new_n240_), .ZN(G1336gat));
  NAND3_X1  g499(.A1(new_n694_), .A2(new_n442_), .A3(new_n376_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n634_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n442_), .ZN(G1337gat));
  OAI21_X1  g502(.A(G99gat), .B1(new_n696_), .B2(new_n356_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n355_), .A2(new_n446_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n693_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g506(.A1(new_n694_), .A2(new_n399_), .A3(new_n370_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n614_), .A2(new_n543_), .A3(new_n370_), .A4(new_n662_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G106gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G106gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT53), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT53), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n708_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1339gat));
  NOR3_X1   g516(.A1(new_n376_), .A2(new_n245_), .A3(new_n379_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n511_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n615_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n502_), .A2(new_n504_), .A3(new_n493_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n509_), .A2(KEYINPUT55), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n505_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n723_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n510_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n502_), .A2(new_n504_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n730_), .B2(new_n492_), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT55), .B(new_n493_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n722_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT56), .B1(new_n733_), .B2(new_n482_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n721_), .B1(new_n729_), .B2(new_n734_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .A4(new_n564_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n553_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n548_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n563_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n506_), .B2(new_n511_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(KEYINPUT115), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n743_), .B(new_n740_), .C1(new_n506_), .C2(new_n511_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n735_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(KEYINPUT57), .A3(new_n625_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n728_), .B1(new_n727_), .B2(new_n510_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n733_), .A2(KEYINPUT56), .A3(new_n482_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n740_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n511_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT58), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n755_), .B(new_n752_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n754_), .A2(new_n756_), .A3(new_n476_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n747_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n750_), .A2(new_n753_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n755_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n750_), .A2(KEYINPUT58), .A3(new_n753_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n758_), .A3(new_n611_), .A4(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n565_), .A2(new_n511_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n741_), .B(KEYINPUT115), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n625_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n763_), .A2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n543_), .B1(new_n759_), .B2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n476_), .A2(new_n615_), .A3(new_n544_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT54), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT54), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n719_), .B1(new_n771_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G113gat), .B1(new_n777_), .B2(new_n565_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT117), .Z(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT57), .B1(new_n746_), .B2(new_n625_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT118), .B1(new_n757_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n761_), .A2(new_n611_), .A3(new_n762_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n769_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n747_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n775_), .B1(new_n786_), .B2(new_n543_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n718_), .A2(new_n780_), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n777_), .A2(new_n780_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n565_), .A2(G113gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n779_), .B1(new_n790_), .B2(new_n791_), .ZN(G1340gat));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n789_), .B2(new_n661_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n786_), .A2(new_n543_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n776_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n788_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n783_), .A2(KEYINPUT116), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n799_), .A2(new_n763_), .A3(new_n769_), .A4(new_n747_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n775_), .B1(new_n800_), .B2(new_n543_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT59), .B1(new_n801_), .B2(new_n719_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n798_), .A2(KEYINPUT119), .A3(new_n516_), .A4(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n794_), .A2(G120gat), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT60), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n661_), .B2(G120gat), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n777_), .B(new_n806_), .C1(new_n805_), .C2(G120gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT120), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(new_n810_), .A3(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1341gat));
  INV_X1    g611(.A(G127gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n789_), .B1(KEYINPUT121), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  OAI21_X1  g614(.A(G127gat), .B1(new_n543_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n777_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n814_), .A2(new_n816_), .B1(new_n813_), .B2(new_n817_), .ZN(G1342gat));
  AOI21_X1  g617(.A(G134gat), .B1(new_n777_), .B2(new_n576_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n611_), .A2(G134gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n790_), .B2(new_n820_), .ZN(G1343gat));
  NOR4_X1   g620(.A1(new_n801_), .A2(new_n245_), .A3(new_n378_), .A4(new_n674_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n565_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT122), .B(G141gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1344gat));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n516_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g626(.A1(new_n822_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT61), .B(G155gat), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1346gat));
  AOI21_X1  g629(.A(G162gat), .B1(new_n822_), .B2(new_n576_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n611_), .A2(G162gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n822_), .B2(new_n832_), .ZN(G1347gat));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n634_), .A2(new_n244_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n355_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n795_), .B2(new_n776_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n260_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n837_), .A2(new_n565_), .A3(new_n371_), .A4(new_n838_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n787_), .A2(new_n615_), .A3(new_n370_), .A4(new_n836_), .ZN(new_n840_));
  INV_X1    g639(.A(G169gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT62), .ZN(new_n843_));
  INV_X1    g642(.A(new_n836_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n796_), .A2(new_n565_), .A3(new_n371_), .A4(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT62), .B1(new_n845_), .B2(G169gat), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n834_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(G169gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n839_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n851_), .A2(KEYINPUT123), .A3(new_n846_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n848_), .A2(new_n852_), .ZN(G1348gat));
  NOR4_X1   g652(.A1(new_n801_), .A2(new_n301_), .A3(new_n661_), .A4(new_n370_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n844_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n787_), .A2(new_n370_), .A3(new_n836_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n856_), .A2(new_n516_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(G176gat), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1349gat));
  OR4_X1    g659(.A1(new_n543_), .A2(new_n801_), .A3(new_n370_), .A4(new_n836_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n543_), .A2(new_n267_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n861_), .A2(new_n293_), .B1(new_n856_), .B2(new_n862_), .ZN(G1350gat));
  NAND3_X1  g662(.A1(new_n856_), .A2(new_n266_), .A3(new_n576_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n856_), .A2(new_n611_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n251_), .ZN(G1351gat));
  NOR2_X1   g665(.A1(new_n801_), .A2(new_n378_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n835_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n615_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT125), .B(G197gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1352gat));
  NOR2_X1   g670(.A1(new_n868_), .A2(new_n661_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n281_), .ZN(G1353gat));
  NOR2_X1   g672(.A1(new_n868_), .A2(new_n543_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT63), .B(G211gat), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n874_), .B2(new_n876_), .ZN(G1354gat));
  XOR2_X1   g676(.A(KEYINPUT126), .B(G218gat), .Z(new_n878_));
  NOR3_X1   g677(.A1(new_n868_), .A2(new_n476_), .A3(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n867_), .A2(new_n576_), .A3(new_n835_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n878_), .ZN(G1355gat));
endmodule


