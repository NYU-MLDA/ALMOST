//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n985_, new_n987_, new_n988_, new_n990_,
    new_n991_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1002_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1009_, new_n1010_, new_n1011_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT5), .B(G176gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT10), .B(G99gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G106gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT65), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n209_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  AND3_X1   g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT9), .A3(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(KEYINPUT9), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n222_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n218_), .A2(new_n219_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n219_), .B1(new_n218_), .B2(new_n229_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(KEYINPUT11), .B2(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n221_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .A4(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n225_), .A2(new_n226_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT8), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n249_), .B1(new_n246_), .B2(KEYINPUT67), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n245_), .A2(KEYINPUT67), .A3(new_n249_), .A4(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n232_), .A2(new_n233_), .A3(new_n238_), .A4(new_n253_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT65), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n216_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n229_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT66), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n218_), .A2(new_n219_), .A3(new_n229_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n238_), .A3(new_n253_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT68), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n258_), .A2(new_n253_), .A3(new_n259_), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n236_), .B(new_n237_), .Z(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT69), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n260_), .A2(new_n266_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n262_), .A2(new_n274_), .A3(new_n263_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n206_), .B1(new_n272_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n265_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n270_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n277_), .B(new_n206_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(KEYINPUT13), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT13), .B1(new_n279_), .B2(new_n282_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT15), .ZN(new_n288_));
  XOR2_X1   g087(.A(G29gat), .B(G36gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(G43gat), .B(G50gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G43gat), .B(G50gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n288_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n294_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n295_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT15), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G1gat), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT77), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(KEYINPUT14), .C1(new_n304_), .C2(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G15gat), .B(G22gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G1gat), .B(G8gat), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n310_), .B(new_n316_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n298_), .A2(new_n303_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n302_), .A4(new_n301_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G229gat), .A2(G233gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n301_), .A2(new_n302_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n322_), .B1(new_n327_), .B2(new_n321_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n287_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n322_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n321_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n318_), .A2(new_n319_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(KEYINPUT79), .C1(new_n320_), .C2(new_n323_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G169gat), .B(G197gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G141gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT80), .B(G113gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n329_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(KEYINPUT81), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n333_), .B(new_n338_), .C1(new_n320_), .C2(new_n323_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT82), .ZN(new_n343_));
  INV_X1    g142(.A(new_n324_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n333_), .A4(new_n338_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n340_), .A2(KEYINPUT81), .B1(new_n343_), .B2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n286_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n325_), .B(new_n263_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G231gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT78), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G127gat), .B(G155gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT16), .ZN(new_n356_));
  INV_X1    g155(.A(G183gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G211gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT17), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n354_), .B(new_n361_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n353_), .A2(KEYINPUT17), .A3(new_n360_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n350_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT87), .ZN(new_n368_));
  XOR2_X1   g167(.A(G71gat), .B(G99gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G15gat), .B(G43gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT24), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(G169gat), .B2(G176gat), .ZN(new_n375_));
  INV_X1    g174(.A(G169gat), .ZN(new_n376_));
  INV_X1    g175(.A(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT85), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT85), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(G183gat), .A3(G190gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT23), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(G183gat), .B2(G190gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n379_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G190gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT26), .B1(new_n389_), .B2(KEYINPUT84), .ZN(new_n390_));
  OR3_X1    g189(.A1(new_n389_), .A2(KEYINPUT84), .A3(KEYINPUT26), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT83), .B(G183gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n390_), .B(new_n391_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n380_), .A2(new_n385_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n381_), .A2(new_n383_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(KEYINPUT23), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n389_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT22), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G169gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n376_), .A2(KEYINPUT22), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT86), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408_));
  AOI21_X1  g207(.A(G176gat), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n407_), .A2(new_n409_), .B1(G169gat), .B2(G176gat), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n388_), .A2(new_n396_), .B1(new_n402_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT30), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n399_), .A2(KEYINPUT23), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n413_), .A2(new_n401_), .A3(new_n397_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n391_), .A2(new_n390_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n357_), .A2(KEYINPUT83), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n357_), .A2(KEYINPUT83), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT25), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n395_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI22_X1  g222(.A1(new_n414_), .A2(new_n417_), .B1(new_n423_), .B2(new_n387_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n412_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n412_), .A3(KEYINPUT88), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n372_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n372_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G127gat), .B(G134gat), .Z(new_n434_));
  XOR2_X1   g233(.A(G113gat), .B(G120gat), .Z(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT31), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n431_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT91), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G155gat), .B(G162gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(KEYINPUT1), .ZN(new_n445_));
  INV_X1    g244(.A(G141gat), .ZN(new_n446_));
  INV_X1    g245(.A(G148gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G141gat), .A2(G148gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT3), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT3), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(G141gat), .B2(G148gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n450_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT2), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT2), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n450_), .B2(new_n460_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n456_), .B(new_n458_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n444_), .B1(new_n464_), .B2(KEYINPUT90), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n450_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT89), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n461_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n453_), .A2(new_n455_), .B1(new_n457_), .B2(KEYINPUT2), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT90), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  AOI211_X1 g270(.A(new_n443_), .B(new_n452_), .C1(new_n465_), .C2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(KEYINPUT90), .ZN(new_n473_));
  INV_X1    g272(.A(new_n444_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n452_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT91), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n442_), .B1(new_n478_), .B2(KEYINPUT29), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G22gat), .B(G50gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n468_), .A2(new_n470_), .A3(new_n469_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n470_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n444_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n443_), .B1(new_n483_), .B2(new_n452_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n475_), .A2(KEYINPUT91), .A3(new_n476_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n487_));
  INV_X1    g286(.A(new_n442_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n479_), .A2(new_n480_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n480_), .B1(new_n479_), .B2(new_n489_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(G228gat), .A2(G233gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n487_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n203_), .B2(G197gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n203_), .A2(G197gat), .ZN(new_n497_));
  INV_X1    g296(.A(G197gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT21), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n203_), .A2(G197gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n498_), .A2(G204gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT21), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G211gat), .B(G218gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n505_), .B(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n500_), .A2(KEYINPUT21), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n501_), .A2(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n493_), .B1(new_n494_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT95), .B(new_n493_), .C1(new_n494_), .C2(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n510_), .A2(new_n493_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT97), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n515_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n492_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n519_), .A2(KEYINPUT96), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(KEYINPUT96), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n515_), .A2(new_n527_), .A3(new_n517_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n526_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n441_), .B(new_n525_), .C1(new_n531_), .C2(new_n492_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G225gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT4), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n484_), .A2(new_n436_), .A3(new_n485_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n483_), .A2(new_n436_), .A3(new_n452_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT4), .B1(new_n478_), .B2(new_n436_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n535_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G1gat), .B(G29gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G57gat), .B(G85gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  NAND3_X1  g346(.A1(new_n537_), .A2(new_n534_), .A3(new_n539_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT102), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT102), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n537_), .A2(new_n550_), .A3(new_n539_), .A4(new_n534_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n542_), .A2(new_n547_), .A3(new_n549_), .A4(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT33), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n549_), .A2(new_n551_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n555_), .A2(KEYINPUT33), .A3(new_n547_), .A4(new_n542_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G8gat), .B(G36gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT18), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G64gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n224_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n404_), .A2(new_n405_), .A3(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n564_), .A3(new_n377_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n416_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n357_), .A2(new_n389_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT100), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT100), .B(new_n567_), .C1(new_n384_), .C2(new_n386_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n566_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT25), .B(G183gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G190gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n400_), .A2(new_n379_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT98), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n400_), .A2(new_n578_), .A3(new_n379_), .A4(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n506_), .A2(new_n501_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n508_), .A2(new_n509_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n572_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G226gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT19), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(KEYINPUT20), .B(new_n587_), .C1(new_n411_), .C2(new_n510_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n583_), .B1(new_n572_), .B2(new_n580_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT20), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n411_), .B2(new_n510_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n587_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n561_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n577_), .A2(new_n579_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n570_), .A2(new_n571_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n566_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n510_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n591_), .B1(new_n424_), .B2(new_n583_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n587_), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT20), .B1(new_n424_), .B2(new_n583_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n595_), .A2(new_n598_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n583_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n601_), .B(new_n560_), .C1(new_n604_), .C2(new_n587_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n594_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n534_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n436_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n472_), .A2(new_n477_), .A3(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n538_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n547_), .B1(new_n610_), .B2(new_n535_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n606_), .B1(new_n607_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n554_), .A2(new_n556_), .A3(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n598_), .A2(new_n510_), .A3(new_n576_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT20), .B1(new_n411_), .B2(new_n510_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n586_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n590_), .A2(new_n592_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n616_), .B1(new_n586_), .B2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n560_), .A2(KEYINPUT32), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n601_), .B1(new_n604_), .B2(new_n587_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n619_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n547_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT4), .B1(new_n609_), .B2(new_n538_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n537_), .A2(new_n536_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n534_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n549_), .A2(new_n551_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n622_), .B1(new_n628_), .B2(new_n552_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n613_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT103), .B(new_n622_), .C1(new_n628_), .C2(new_n552_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n533_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n525_), .B1(new_n531_), .B2(new_n492_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n441_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n618_), .A2(new_n561_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT27), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n589_), .A2(new_n593_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n560_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n637_), .A2(new_n640_), .B1(new_n606_), .B2(new_n638_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n628_), .A3(new_n552_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n532_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n633_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n298_), .A2(new_n303_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n262_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT74), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n296_), .A2(new_n297_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n649_), .A2(new_n258_), .A3(new_n253_), .A4(new_n259_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT34), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT35), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .A4(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT72), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT72), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n647_), .A2(new_n658_), .A3(new_n650_), .A4(new_n655_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n653_), .A2(new_n654_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n647_), .A2(new_n650_), .A3(new_n655_), .ZN(new_n662_));
  OAI221_X1 g461(.A(KEYINPUT72), .B1(new_n654_), .B2(new_n653_), .C1(new_n662_), .C2(KEYINPUT74), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(G190gat), .B(G218gat), .Z(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT73), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(G134gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(G162gat), .Z(new_n668_));
  INV_X1    g467(.A(KEYINPUT36), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n664_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT37), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n669_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n664_), .A2(KEYINPUT75), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT75), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n663_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n670_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n674_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n675_), .B1(new_n682_), .B2(new_n672_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n366_), .A2(new_n645_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT104), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n628_), .A2(new_n552_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n622_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT103), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n629_), .A2(new_n630_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n613_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n530_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n692_), .A2(new_n528_), .B1(KEYINPUT96), .B2(new_n519_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n492_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n523_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n693_), .A2(new_n694_), .B1(new_n695_), .B2(new_n522_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n642_), .B1(new_n696_), .B2(new_n441_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n691_), .A2(new_n533_), .B1(new_n636_), .B2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n698_), .A2(new_n350_), .A3(new_n365_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n683_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n685_), .A2(new_n701_), .A3(new_n304_), .A4(new_n686_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT38), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(new_n686_), .A3(new_n682_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G1gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n703_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n706_), .A3(new_n707_), .ZN(G1324gat));
  INV_X1    g507(.A(new_n641_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n366_), .A2(new_n709_), .A3(new_n645_), .A4(new_n682_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G8gat), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT39), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT105), .B1(new_n710_), .B2(G8gat), .ZN(new_n715_));
  OR3_X1    g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n685_), .A2(new_n701_), .A3(new_n305_), .A4(new_n709_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n714_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n716_), .A2(KEYINPUT40), .A3(new_n717_), .A4(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n717_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n719_), .A2(new_n723_), .ZN(G1325gat));
  INV_X1    g523(.A(new_n684_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n441_), .A2(G15gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(KEYINPUT106), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728_));
  INV_X1    g527(.A(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n684_), .B2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n727_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n699_), .A2(new_n635_), .A3(new_n682_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G15gat), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n732_), .A3(G15gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT107), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n731_), .A2(new_n739_), .A3(new_n735_), .A4(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1326gat));
  OR3_X1    g540(.A1(new_n684_), .A2(G22gat), .A3(new_n696_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n699_), .A2(new_n634_), .A3(new_n682_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G22gat), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT108), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(KEYINPUT108), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(KEYINPUT42), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT42), .B1(new_n745_), .B2(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n742_), .B1(new_n747_), .B2(new_n748_), .ZN(G1327gat));
  NOR2_X1   g548(.A1(new_n350_), .A2(new_n364_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n670_), .B1(new_n664_), .B2(KEYINPUT75), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n674_), .B1(new_n752_), .B2(new_n678_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n681_), .A2(KEYINPUT37), .ZN(new_n754_));
  OAI22_X1  g553(.A1(new_n753_), .A2(KEYINPUT37), .B1(new_n671_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n645_), .B2(new_n755_), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT43), .B(new_n683_), .C1(new_n633_), .C2(new_n644_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT44), .B(new_n750_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(G29gat), .A3(new_n686_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT43), .B1(new_n698_), .B2(new_n683_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n645_), .A2(new_n751_), .A3(new_n755_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT44), .B1(new_n762_), .B2(new_n750_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n698_), .A2(new_n682_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n750_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n686_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n759_), .A2(new_n763_), .B1(G29gat), .B2(new_n767_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT109), .Z(G1328gat));
  NAND2_X1  g568(.A1(new_n758_), .A2(new_n709_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G36gat), .B1(new_n770_), .B2(new_n763_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n641_), .A2(G36gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n750_), .A3(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT110), .B(KEYINPUT112), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n764_), .A2(new_n750_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n778_));
  AND3_X1   g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n771_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n771_), .B(KEYINPUT46), .C1(new_n779_), .C2(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1329gat));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  INV_X1    g586(.A(G43gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n765_), .B2(new_n441_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n441_), .A2(new_n788_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n758_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n787_), .B(new_n789_), .C1(new_n791_), .C2(new_n763_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n750_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n758_), .A3(new_n790_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n787_), .B1(new_n797_), .B2(new_n789_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n786_), .B1(new_n793_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n789_), .B1(new_n791_), .B2(new_n763_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT113), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT47), .A3(new_n792_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(G1330gat));
  INV_X1    g602(.A(new_n765_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G50gat), .B1(new_n804_), .B2(new_n634_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n758_), .A2(G50gat), .A3(new_n634_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n796_), .ZN(G1331gat));
  NAND2_X1  g606(.A1(new_n364_), .A2(new_n348_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n698_), .A2(new_n286_), .A3(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n682_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(G57gat), .A3(new_n686_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(G57gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n809_), .A2(new_n683_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n766_), .B1(new_n815_), .B2(KEYINPUT114), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(KEYINPUT114), .B2(new_n815_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n814_), .B2(new_n817_), .ZN(G1332gat));
  INV_X1    g617(.A(G64gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n810_), .B2(new_n709_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT48), .Z(new_n821_));
  INV_X1    g620(.A(new_n815_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n819_), .A3(new_n709_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1333gat));
  INV_X1    g623(.A(G71gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n810_), .B2(new_n635_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT49), .Z(new_n827_));
  NAND3_X1  g626(.A1(new_n822_), .A2(new_n825_), .A3(new_n635_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1334gat));
  OR3_X1    g628(.A1(new_n815_), .A2(G78gat), .A3(new_n696_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n810_), .A2(new_n634_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G78gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n833_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n830_), .B1(new_n834_), .B2(new_n835_), .ZN(G1335gat));
  NOR3_X1   g635(.A1(new_n286_), .A2(new_n364_), .A3(new_n349_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n764_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n223_), .A3(new_n686_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n762_), .A2(new_n837_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n840_), .A2(new_n686_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n841_), .B2(new_n223_), .ZN(G1336gat));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n224_), .A3(new_n709_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n840_), .A2(new_n709_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n224_), .ZN(G1337gat));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n635_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G99gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n838_), .A2(new_n635_), .A3(new_n212_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT51), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n851_), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1338gat));
  NAND3_X1  g652(.A1(new_n838_), .A2(new_n634_), .A3(new_n215_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n762_), .A2(new_n634_), .A3(new_n837_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(G106gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n855_), .B2(G106gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT118), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n854_), .B(new_n861_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1339gat));
  NOR3_X1   g664(.A1(new_n766_), .A2(new_n709_), .A3(new_n441_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n277_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n273_), .B(KEYINPUT55), .C1(new_n275_), .C2(new_n276_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n261_), .B(new_n254_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n267_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(KEYINPUT119), .A3(new_n267_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n870_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI22_X1  g675(.A1(new_n876_), .A2(new_n206_), .B1(KEYINPUT120), .B2(KEYINPUT56), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n871_), .A2(KEYINPUT119), .A3(new_n267_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT119), .B1(new_n871_), .B2(new_n267_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n868_), .B(new_n869_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n206_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n275_), .A2(new_n276_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n269_), .A2(new_n271_), .B1(new_n884_), .B2(new_n273_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n341_), .A2(new_n347_), .B1(new_n885_), .B2(new_n206_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n877_), .A2(new_n883_), .A3(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n320_), .A2(new_n331_), .A3(new_n322_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n322_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n339_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n890_), .B2(KEYINPUT121), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n890_), .A2(KEYINPUT121), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n891_), .A2(new_n892_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n282_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n278_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n893_), .B(KEYINPUT122), .C1(new_n278_), .C2(new_n894_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n887_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n899_), .A2(KEYINPUT57), .A3(new_n682_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n899_), .B2(new_n682_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n876_), .B2(new_n206_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n880_), .A2(KEYINPUT56), .A3(new_n881_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n893_), .A2(new_n282_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT58), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n903_), .B1(new_n910_), .B2(new_n683_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n755_), .B(KEYINPUT123), .C1(new_n912_), .C2(KEYINPUT58), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(KEYINPUT58), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n364_), .B1(new_n902_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n285_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n283_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n808_), .ZN(new_n919_));
  AOI21_X1  g718(.A(KEYINPUT54), .B1(new_n919_), .B2(new_n683_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n918_), .A2(new_n755_), .A3(new_n921_), .A4(new_n808_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n920_), .A2(new_n922_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n696_), .B(new_n866_), .C1(new_n916_), .C2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT59), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n899_), .A2(new_n682_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n899_), .A2(KEYINPUT57), .A3(new_n682_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n365_), .B1(new_n926_), .B2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n920_), .A2(new_n922_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT59), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n934_), .A2(new_n935_), .A3(new_n696_), .A4(new_n866_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n925_), .A2(new_n936_), .A3(new_n349_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G113gat), .ZN(new_n938_));
  OR3_X1    g737(.A1(new_n924_), .A2(G113gat), .A3(new_n348_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1340gat));
  NAND3_X1  g739(.A1(new_n925_), .A2(new_n936_), .A3(new_n918_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(G120gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n634_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(G120gat), .ZN(new_n945_));
  AOI21_X1  g744(.A(G120gat), .B1(new_n918_), .B2(new_n944_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(KEYINPUT124), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(KEYINPUT124), .B2(new_n946_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n943_), .A2(new_n866_), .A3(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n942_), .A2(new_n949_), .ZN(G1341gat));
  NAND3_X1  g749(.A1(new_n925_), .A2(new_n936_), .A3(new_n364_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(G127gat), .ZN(new_n952_));
  OR3_X1    g751(.A1(new_n924_), .A2(G127gat), .A3(new_n365_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1342gat));
  NAND3_X1  g753(.A1(new_n925_), .A2(new_n936_), .A3(new_n755_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(G134gat), .ZN(new_n956_));
  OR3_X1    g755(.A1(new_n924_), .A2(G134gat), .A3(new_n682_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1343gat));
  NOR2_X1   g757(.A1(new_n696_), .A2(new_n635_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n960_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n766_), .A2(new_n709_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n961_), .A2(new_n349_), .A3(new_n962_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g763(.A1(new_n961_), .A2(new_n918_), .A3(new_n962_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g765(.A1(new_n961_), .A2(new_n364_), .A3(new_n962_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(KEYINPUT61), .B(G155gat), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(KEYINPUT125), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n967_), .B(new_n969_), .ZN(G1346gat));
  NAND2_X1  g769(.A1(new_n961_), .A2(new_n962_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G162gat), .B1(new_n971_), .B2(new_n683_), .ZN(new_n972_));
  OR2_X1    g771(.A1(new_n682_), .A2(G162gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n971_), .B2(new_n973_), .ZN(G1347gat));
  NOR3_X1   g773(.A1(new_n686_), .A2(new_n441_), .A3(new_n641_), .ZN(new_n975_));
  OAI211_X1 g774(.A(new_n696_), .B(new_n975_), .C1(new_n916_), .C2(new_n923_), .ZN(new_n976_));
  OAI21_X1  g775(.A(G169gat), .B1(new_n976_), .B2(new_n348_), .ZN(new_n977_));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n977_), .A2(new_n978_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n943_), .A2(new_n349_), .A3(new_n975_), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n980_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n981_));
  AND2_X1   g780(.A1(new_n562_), .A2(new_n564_), .ZN(new_n982_));
  INV_X1    g781(.A(new_n982_), .ZN(new_n983_));
  OAI211_X1 g782(.A(new_n979_), .B(new_n981_), .C1(new_n980_), .C2(new_n983_), .ZN(G1348gat));
  NOR2_X1   g783(.A1(new_n976_), .A2(new_n286_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(new_n377_), .ZN(G1349gat));
  NAND3_X1  g785(.A1(new_n943_), .A2(new_n364_), .A3(new_n975_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(new_n987_), .A2(new_n573_), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n988_), .B1(new_n392_), .B2(new_n987_), .ZN(G1350gat));
  OAI21_X1  g788(.A(G190gat), .B1(new_n976_), .B2(new_n683_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n753_), .A2(new_n574_), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n990_), .B1(new_n976_), .B2(new_n991_), .ZN(G1351gat));
  NOR2_X1   g791(.A1(new_n686_), .A2(new_n641_), .ZN(new_n993_));
  NAND4_X1  g792(.A1(new_n961_), .A2(G197gat), .A3(new_n349_), .A4(new_n993_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n994_), .A2(KEYINPUT126), .ZN(new_n995_));
  OAI211_X1 g794(.A(new_n959_), .B(new_n993_), .C1(new_n916_), .C2(new_n923_), .ZN(new_n996_));
  INV_X1    g795(.A(new_n996_), .ZN(new_n997_));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n998_));
  NAND4_X1  g797(.A1(new_n997_), .A2(new_n998_), .A3(G197gat), .A4(new_n349_), .ZN(new_n999_));
  OAI21_X1  g798(.A(new_n498_), .B1(new_n996_), .B2(new_n348_), .ZN(new_n1000_));
  AND3_X1   g799(.A1(new_n995_), .A2(new_n999_), .A3(new_n1000_), .ZN(G1352gat));
  NOR2_X1   g800(.A1(new_n996_), .A2(new_n286_), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(new_n1002_), .B(new_n203_), .ZN(G1353gat));
  NOR2_X1   g802(.A1(new_n996_), .A2(new_n365_), .ZN(new_n1004_));
  NOR2_X1   g803(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1005_));
  AND2_X1   g804(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1006_));
  OAI21_X1  g805(.A(new_n1004_), .B1(new_n1005_), .B2(new_n1006_), .ZN(new_n1007_));
  OAI21_X1  g806(.A(new_n1007_), .B1(new_n1004_), .B2(new_n1005_), .ZN(G1354gat));
  AOI21_X1  g807(.A(G218gat), .B1(new_n997_), .B2(new_n753_), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n755_), .A2(G218gat), .ZN(new_n1010_));
  XNOR2_X1  g809(.A(new_n1010_), .B(KEYINPUT127), .ZN(new_n1011_));
  AOI21_X1  g810(.A(new_n1009_), .B1(new_n997_), .B2(new_n1011_), .ZN(G1355gat));
endmodule


