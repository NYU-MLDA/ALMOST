//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT79), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT79), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT24), .A4(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT26), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G190gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n215_), .A2(new_n217_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n202_), .A3(new_n203_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n208_), .A2(new_n213_), .A3(new_n222_), .A4(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n211_), .B(new_n212_), .C1(G183gat), .C2(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n202_), .A2(KEYINPUT22), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G169gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n229_), .A3(new_n203_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n207_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT87), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT21), .B(new_n233_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  INV_X1    g036(.A(G218gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G211gat), .ZN(new_n239_));
  INV_X1    g038(.A(G211gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G218gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n237_), .B1(new_n242_), .B2(KEYINPUT87), .ZN(new_n243_));
  AND2_X1   g042(.A1(G197gat), .A2(G204gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G197gat), .A2(G204gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n234_), .B2(KEYINPUT21), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n236_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n232_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT19), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(KEYINPUT88), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n230_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n227_), .A2(new_n229_), .A3(KEYINPUT80), .A4(new_n203_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n255_), .A2(new_n226_), .A3(new_n207_), .A4(new_n256_), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n205_), .A2(G169gat), .A3(G176gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT79), .B1(new_n202_), .B2(new_n203_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n223_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n260_), .A2(new_n213_), .A3(new_n208_), .A4(new_n222_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n263_), .B(new_n236_), .C1(new_n243_), .C2(new_n247_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT20), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n252_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n262_), .B1(new_n253_), .B2(new_n264_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n257_), .A2(new_n261_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n264_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n240_), .A2(G218gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n238_), .A2(G211gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n237_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n235_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n276_), .B(new_n246_), .C1(new_n277_), .C2(new_n237_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n263_), .B1(new_n278_), .B2(new_n236_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n272_), .B1(new_n273_), .B2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n232_), .A2(new_n248_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n271_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n267_), .B1(new_n283_), .B2(new_n251_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT18), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT94), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n284_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n284_), .A2(KEYINPUT94), .A3(new_n288_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT89), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n248_), .B(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(new_n232_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n251_), .B1(new_n301_), .B2(new_n266_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n283_), .B2(new_n251_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n293_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(new_n289_), .A3(KEYINPUT27), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT3), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT2), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(KEYINPUT1), .B2(new_n312_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(KEYINPUT1), .B2(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n309_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(new_n307_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n311_), .A2(new_n315_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT85), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n311_), .A2(new_n315_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n317_), .A2(new_n319_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT28), .B1(new_n329_), .B2(KEYINPUT29), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G22gat), .B(G50gat), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n300_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT90), .Z(new_n345_));
  XOR2_X1   g144(.A(new_n341_), .B(KEYINPUT86), .Z(new_n346_));
  NAND4_X1  g145(.A1(new_n339_), .A2(new_n264_), .A3(new_n253_), .A4(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n343_), .A2(KEYINPUT91), .A3(new_n345_), .A4(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n343_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT91), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n338_), .B(new_n348_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n326_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n334_), .B1(new_n326_), .B2(new_n332_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT92), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n349_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n343_), .A2(new_n347_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n344_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n343_), .A2(KEYINPUT92), .A3(new_n345_), .A4(new_n347_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n356_), .A2(new_n358_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n353_), .A2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n306_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT81), .B(G43gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n272_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(G15gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT30), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n368_), .B(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT83), .ZN(new_n374_));
  XOR2_X1   g173(.A(G127gat), .B(G134gat), .Z(new_n375_));
  XOR2_X1   g174(.A(G113gat), .B(G120gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT82), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n373_), .A2(KEYINPUT83), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n382_), .A3(new_n380_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT95), .ZN(new_n385_));
  INV_X1    g184(.A(new_n377_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n329_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n329_), .A2(new_n386_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n320_), .A2(new_n377_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(KEYINPUT4), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n385_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G1gat), .B(G29gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT96), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT0), .B(G57gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n393_), .A3(new_n389_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n394_), .A2(new_n385_), .A3(new_n390_), .A4(new_n388_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n396_), .A2(new_n402_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n403_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n401_), .B1(new_n406_), .B2(new_n395_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n384_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n364_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n284_), .A2(KEYINPUT94), .A3(new_n288_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT94), .B1(new_n284_), .B2(new_n288_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n284_), .A2(new_n288_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n412_), .B(new_n305_), .C1(new_n416_), .C2(KEYINPUT27), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT100), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n298_), .A2(KEYINPUT100), .A3(new_n412_), .A4(new_n305_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n288_), .A2(KEYINPUT32), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n303_), .A2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n408_), .B(new_n422_), .C1(new_n292_), .C2(new_n421_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n405_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n406_), .A2(new_n395_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(KEYINPUT33), .A3(new_n402_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n394_), .A2(new_n389_), .A3(new_n388_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT98), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n394_), .A2(KEYINPUT98), .A3(new_n389_), .A4(new_n388_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n392_), .A2(new_n393_), .A3(new_n390_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n401_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(KEYINPUT97), .A3(new_n401_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n432_), .A2(new_n438_), .A3(KEYINPUT99), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT99), .B1(new_n432_), .B2(new_n438_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n425_), .B(new_n427_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n423_), .B1(new_n441_), .B2(new_n296_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n363_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n419_), .A2(new_n420_), .A3(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n384_), .B(KEYINPUT84), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT101), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n411_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G15gat), .B(G22gat), .ZN(new_n452_));
  INV_X1    g251(.A(G1gat), .ZN(new_n453_));
  INV_X1    g252(.A(G8gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT14), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G1gat), .B(G8gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  XOR2_X1   g257(.A(G29gat), .B(G36gat), .Z(new_n459_));
  XOR2_X1   g258(.A(G43gat), .B(G50gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n456_), .B(new_n457_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G229gat), .A2(G233gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n465_), .A3(KEYINPUT76), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n461_), .B(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n464_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n469_), .A3(new_n462_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT77), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT78), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT78), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(KEYINPUT77), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G169gat), .B(G197gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n484_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n480_), .B1(new_n477_), .B2(KEYINPUT77), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT77), .ZN(new_n488_));
  AOI211_X1 g287(.A(new_n488_), .B(KEYINPUT78), .C1(new_n472_), .C2(new_n476_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G190gat), .B(G218gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G134gat), .B(G162gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(KEYINPUT36), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(KEYINPUT35), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT64), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n504_), .B(KEYINPUT7), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT64), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G85gat), .B(G92gat), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT8), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n512_), .B1(new_n506_), .B2(new_n503_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT10), .B(G99gat), .Z(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  AOI22_X1  g318(.A1(KEYINPUT9), .A2(new_n512_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT9), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n503_), .A2(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n516_), .A2(new_n517_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n515_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n500_), .B1(new_n474_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n517_), .A2(new_n516_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n513_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n461_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n499_), .A2(KEYINPUT35), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT68), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n536_), .A2(new_n537_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n527_), .A2(new_n537_), .A3(new_n536_), .A4(new_n533_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n497_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n540_), .A2(new_n497_), .A3(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n495_), .A2(KEYINPUT36), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT72), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT37), .B1(new_n542_), .B2(KEYINPUT71), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n551_));
  INV_X1    g350(.A(new_n544_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n551_), .B(new_n546_), .C1(new_n552_), .C2(new_n542_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n549_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT74), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G127gat), .B(G155gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n464_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT65), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(KEYINPUT11), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n573_));
  XOR2_X1   g372(.A(G71gat), .B(G78gat), .Z(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n569_), .A3(KEYINPUT11), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(KEYINPUT11), .B2(new_n570_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n578_), .B2(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n568_), .B(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n566_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n564_), .A2(new_n565_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n566_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT75), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n558_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n532_), .A2(new_n580_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n580_), .A2(new_n515_), .A3(new_n525_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n589_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n532_), .B2(new_n580_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n580_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n526_), .A2(KEYINPUT12), .A3(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n591_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n593_), .B1(new_n598_), .B2(new_n589_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G120gat), .B(G148gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n599_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(KEYINPUT67), .A2(KEYINPUT13), .ZN(new_n606_));
  NOR2_X1   g405(.A1(KEYINPUT67), .A2(KEYINPUT13), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n605_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(KEYINPUT67), .B2(KEYINPUT13), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n587_), .A2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n451_), .A2(new_n492_), .A3(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n408_), .B(KEYINPUT102), .Z(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n453_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n451_), .A2(new_n547_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n610_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n618_), .A2(new_n492_), .A3(new_n585_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n408_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n614_), .A2(new_n615_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n616_), .A2(new_n622_), .A3(new_n623_), .ZN(G1324gat));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n625_));
  INV_X1    g424(.A(new_n306_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G8gat), .B1(new_n620_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n612_), .A2(new_n454_), .A3(new_n306_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT103), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n625_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n627_), .B(KEYINPUT39), .ZN(new_n633_));
  INV_X1    g432(.A(new_n631_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(KEYINPUT40), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n620_), .B2(new_n446_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n446_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n612_), .A2(new_n370_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(G1326gat));
  XNOR2_X1  g442(.A(new_n363_), .B(KEYINPUT105), .ZN(new_n644_));
  OAI21_X1  g443(.A(G22gat), .B1(new_n620_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n644_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n612_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1327gat));
  NOR2_X1   g449(.A1(new_n451_), .A2(new_n492_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n586_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n547_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n618_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n655_), .A2(G29gat), .A3(new_n621_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n558_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT43), .B1(new_n451_), .B2(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n445_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n449_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n410_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n558_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n658_), .A2(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n618_), .A2(new_n492_), .A3(new_n652_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(KEYINPUT44), .A3(new_n665_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n613_), .A3(new_n669_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n670_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT106), .B1(new_n670_), .B2(G29gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n656_), .B1(new_n671_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT44), .B1(new_n664_), .B2(new_n665_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n665_), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n667_), .B(new_n677_), .C1(new_n658_), .C2(new_n663_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n675_), .B1(new_n679_), .B2(new_n306_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n651_), .A2(new_n675_), .A3(new_n306_), .A4(new_n654_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT45), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n674_), .B1(new_n680_), .B2(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n676_), .A2(new_n678_), .A3(new_n626_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT46), .B(new_n682_), .C1(new_n685_), .C2(new_n675_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1329gat));
  INV_X1    g486(.A(G43gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n384_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n668_), .A2(new_n669_), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n655_), .B2(new_n446_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT47), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n690_), .A2(new_n694_), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1330gat));
  NAND2_X1  g495(.A1(new_n679_), .A2(new_n363_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G50gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n644_), .A2(G50gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT107), .Z(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n655_), .B2(new_n700_), .ZN(G1331gat));
  NOR2_X1   g500(.A1(new_n451_), .A2(new_n491_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(new_n618_), .A3(new_n587_), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n613_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n610_), .A2(new_n491_), .A3(new_n586_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n617_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n621_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g508(.A(G64gat), .B1(new_n707_), .B2(new_n626_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n703_), .A2(new_n713_), .A3(new_n306_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n707_), .B2(new_n446_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n446_), .A2(G71gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT109), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n703_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1334gat));
  INV_X1    g520(.A(G78gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n703_), .A2(new_n722_), .A3(new_n648_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G78gat), .B1(new_n707_), .B2(new_n644_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT50), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT50), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT110), .B(new_n723_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n652_), .A2(new_n610_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n653_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n702_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n613_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n521_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT111), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(KEYINPUT111), .ZN(new_n739_));
  INV_X1    g538(.A(new_n664_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n733_), .A2(new_n491_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n621_), .A2(new_n521_), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n738_), .A2(new_n739_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  NOR3_X1   g544(.A1(new_n735_), .A2(G92gat), .A3(new_n626_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n740_), .A2(new_n626_), .A3(new_n742_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n522_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT112), .B(new_n747_), .C1(new_n748_), .C2(new_n522_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1337gat));
  INV_X1    g552(.A(new_n518_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n735_), .A2(new_n384_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n740_), .A2(new_n446_), .A3(new_n742_), .ZN(new_n757_));
  INV_X1    g556(.A(G99gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT51), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n756_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1338gat));
  NAND4_X1  g562(.A1(new_n702_), .A2(new_n519_), .A3(new_n363_), .A4(new_n734_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n664_), .A2(new_n363_), .A3(new_n741_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT53), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n764_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT59), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n599_), .A2(new_n603_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n589_), .B2(KEYINPUT114), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n576_), .A2(new_n579_), .A3(KEYINPUT12), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n591_), .B1(new_n532_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n594_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n526_), .B2(new_n596_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n778_), .B1(new_n777_), .B2(new_n589_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n595_), .A2(new_n591_), .A3(new_n597_), .A4(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT115), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n783_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n603_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n783_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n788_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT56), .B(new_n603_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n491_), .B(new_n776_), .C1(new_n791_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n475_), .A2(new_n470_), .A3(new_n462_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n486_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n477_), .A2(new_n484_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n796_), .A2(new_n797_), .B1(new_n604_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n790_), .A2(new_n603_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n775_), .B1(new_n806_), .B2(new_n794_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT116), .A3(new_n491_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  AND4_X1   g608(.A1(KEYINPUT119), .A2(new_n809_), .A3(KEYINPUT57), .A4(new_n653_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n547_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT119), .B1(new_n811_), .B2(KEYINPUT57), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n653_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n776_), .B(new_n802_), .C1(new_n791_), .C2(new_n795_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n819_), .A2(KEYINPUT58), .B1(new_n554_), .B2(new_n557_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n818_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(KEYINPUT58), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n558_), .A3(new_n823_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT118), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n816_), .A2(new_n824_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n585_), .B1(new_n813_), .B2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n611_), .B2(new_n491_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n587_), .A2(new_n492_), .A3(new_n610_), .A4(new_n830_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n829_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n736_), .A2(new_n384_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n364_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n774_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n838_), .A2(KEYINPUT120), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(KEYINPUT120), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n774_), .A3(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n809_), .A2(KEYINPUT57), .A3(new_n653_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n811_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n816_), .A2(KEYINPUT121), .A3(new_n826_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n811_), .A2(KEYINPUT57), .ZN(new_n851_));
  INV_X1    g650(.A(new_n826_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n849_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n586_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n843_), .B1(new_n855_), .B2(new_n835_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT122), .B1(new_n840_), .B2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n826_), .A2(KEYINPUT118), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n821_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n848_), .A2(new_n860_), .A3(new_n816_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n834_), .B1(new_n861_), .B2(new_n585_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT59), .B1(new_n862_), .B2(new_n838_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  INV_X1    g663(.A(new_n843_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n814_), .A2(new_n815_), .B1(new_n823_), .B2(new_n820_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n866_), .A2(KEYINPUT121), .B1(new_n846_), .B2(new_n847_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n652_), .B1(new_n867_), .B2(new_n853_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n865_), .B1(new_n868_), .B2(new_n834_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n863_), .A2(new_n864_), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n857_), .A2(new_n870_), .A3(new_n491_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G113gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n862_), .A2(new_n838_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OR3_X1    g673(.A1(new_n874_), .A2(G113gat), .A3(new_n492_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(G1340gat));
  XOR2_X1   g675(.A(KEYINPUT123), .B(G120gat), .Z(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n873_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n840_), .A2(new_n856_), .A3(new_n610_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n877_), .ZN(G1341gat));
  INV_X1    g680(.A(new_n585_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n857_), .A2(new_n870_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G127gat), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n874_), .A2(G127gat), .A3(new_n586_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1342gat));
  NAND3_X1  g685(.A1(new_n857_), .A2(new_n870_), .A3(new_n558_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G134gat), .ZN(new_n888_));
  OR3_X1    g687(.A1(new_n874_), .A2(G134gat), .A3(new_n653_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1343gat));
  NOR4_X1   g689(.A1(new_n641_), .A2(new_n443_), .A3(new_n306_), .A4(new_n736_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n836_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n491_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n618_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n892_), .A2(new_n586_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OR3_X1    g699(.A1(new_n892_), .A2(G162gat), .A3(new_n653_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G162gat), .B1(new_n892_), .B2(new_n657_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1347gat));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n834_), .B1(new_n854_), .B2(new_n586_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n446_), .A2(new_n626_), .A3(new_n613_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n644_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n492_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n905_), .A2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n904_), .B1(new_n910_), .B2(new_n202_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT62), .B(G169gat), .C1(new_n905_), .C2(new_n909_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n911_), .A2(new_n912_), .A3(KEYINPUT124), .A4(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1348gat));
  NOR2_X1   g717(.A1(new_n905_), .A2(new_n907_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G176gat), .B1(new_n919_), .B2(new_n618_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n862_), .A2(new_n363_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n906_), .A2(G176gat), .A3(new_n618_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n921_), .A2(new_n652_), .A3(new_n906_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n585_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n924_), .A2(new_n214_), .B1(new_n919_), .B2(new_n925_), .ZN(G1350gat));
  NAND4_X1  g725(.A1(new_n919_), .A2(new_n219_), .A3(new_n221_), .A4(new_n547_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n905_), .A2(new_n657_), .A3(new_n907_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n928_), .B2(new_n218_), .ZN(G1351gat));
  AND3_X1   g728(.A1(new_n446_), .A2(new_n412_), .A3(new_n306_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n836_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n491_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n618_), .ZN(new_n934_));
  INV_X1    g733(.A(G204gat), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(KEYINPUT125), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n934_), .B(new_n936_), .ZN(G1353gat));
  NAND2_X1  g736(.A1(new_n931_), .A2(new_n882_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n941_), .B1(new_n938_), .B2(new_n939_), .ZN(G1354gat));
  AND3_X1   g741(.A1(new_n836_), .A2(new_n547_), .A3(new_n930_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n943_), .A2(KEYINPUT126), .ZN(new_n944_));
  AOI21_X1  g743(.A(G218gat), .B1(new_n943_), .B2(KEYINPUT126), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n657_), .A2(new_n238_), .ZN(new_n946_));
  AOI22_X1  g745(.A1(new_n944_), .A2(new_n945_), .B1(new_n931_), .B2(new_n946_), .ZN(G1355gat));
endmodule


