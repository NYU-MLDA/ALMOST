//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT96), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT91), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT91), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G204gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(G197gat), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT92), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT90), .B(G197gat), .ZN(new_n212_));
  OAI22_X1  g011(.A1(new_n210_), .A2(new_n211_), .B1(G204gat), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT91), .B(G204gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n214_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT21), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT93), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n209_), .A3(new_n217_), .A4(G197gat), .ZN(new_n218_));
  INV_X1    g017(.A(G197gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT90), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G197gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n222_), .A3(G204gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT21), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n207_), .A2(new_n209_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT93), .B1(new_n226_), .B2(new_n219_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n216_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n229_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT21), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  OR3_X1    g039(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT79), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(KEYINPUT79), .A3(new_n241_), .ZN(new_n245_));
  INV_X1    g044(.A(G183gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT25), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G183gat), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT77), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G190gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT26), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(new_n252_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT78), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G169gat), .A3(G176gat), .ZN(new_n262_));
  INV_X1    g061(.A(G169gat), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n262_), .A3(new_n265_), .A4(KEYINPUT24), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n244_), .A2(new_n245_), .A3(new_n258_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(KEYINPUT22), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G169gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n270_), .A3(new_n264_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n260_), .A2(new_n262_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(new_n236_), .B2(KEYINPUT23), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n240_), .B2(new_n273_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n254_), .A2(new_n256_), .A3(new_n246_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n271_), .B(new_n272_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n267_), .A2(KEYINPUT81), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT81), .B1(new_n267_), .B2(new_n277_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n235_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT97), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT80), .B1(new_n237_), .B2(new_n239_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n281_), .B(new_n241_), .C1(new_n282_), .C2(new_n274_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n253_), .A2(KEYINPUT26), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n252_), .A2(new_n247_), .A3(new_n249_), .A4(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n241_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT97), .B1(new_n275_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT98), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n272_), .A2(new_n291_), .A3(new_n271_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n272_), .B2(new_n271_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n246_), .A2(new_n253_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n240_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n295_), .B1(new_n240_), .B2(new_n296_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n288_), .A2(new_n290_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT92), .B1(new_n214_), .B2(G197gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n226_), .A2(new_n211_), .A3(new_n219_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n220_), .A2(new_n222_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n206_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n231_), .B1(new_n305_), .B2(KEYINPUT21), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n233_), .B1(new_n306_), .B2(new_n228_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT20), .B1(new_n300_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n205_), .B1(new_n280_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT20), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(new_n300_), .B2(new_n307_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n235_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n204_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G8gat), .B(G36gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT18), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(new_n314_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT100), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n309_), .A2(KEYINPUT100), .A3(new_n314_), .A4(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n309_), .A2(new_n314_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n318_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT27), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT104), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(KEYINPUT104), .A3(new_n327_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334_));
  OAI22_X1  g133(.A1(new_n333_), .A2(new_n334_), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n334_), .A3(new_n333_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n333_), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n341_), .A2(new_n337_), .A3(KEYINPUT2), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT84), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n341_), .A2(new_n337_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT87), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n352_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT85), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(G141gat), .B2(G148gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n360_));
  AND2_X1   g159(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n357_), .B(new_n359_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n349_), .B1(new_n355_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G127gat), .B(G134gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G113gat), .B(G120gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n347_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n345_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n363_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(new_n371_), .A3(KEYINPUT4), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n369_), .B(new_n373_), .C1(new_n370_), .C2(new_n363_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT101), .B1(new_n372_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n368_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n368_), .A2(new_n371_), .A3(KEYINPUT4), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT101), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n376_), .A4(new_n374_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n378_), .A2(new_n387_), .A3(new_n382_), .A4(new_n379_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n293_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n272_), .A2(new_n291_), .A3(new_n271_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n299_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n290_), .A2(new_n283_), .A3(new_n287_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n310_), .B1(new_n235_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n279_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n267_), .A2(KEYINPUT81), .A3(new_n277_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n307_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n205_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n397_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n313_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n324_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n404_), .A2(KEYINPUT27), .A3(new_n319_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT95), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(KEYINPUT89), .Z(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT29), .B1(new_n370_), .B2(new_n363_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n235_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(KEYINPUT88), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n412_), .B(KEYINPUT29), .C1(new_n370_), .C2(new_n363_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n235_), .A2(new_n411_), .A3(new_n408_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT94), .ZN(new_n415_));
  INV_X1    g214(.A(new_n408_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n230_), .B2(new_n234_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT94), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n410_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n406_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n370_), .A2(new_n363_), .A3(KEYINPUT29), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G22gat), .B(G50gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT28), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n424_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n420_), .A2(new_n422_), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n410_), .B(new_n421_), .C1(new_n415_), .C2(new_n419_), .ZN(new_n430_));
  OAI22_X1  g229(.A1(new_n423_), .A2(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n415_), .A2(new_n419_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n410_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n421_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n420_), .A2(new_n422_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n435_), .A2(new_n406_), .A3(new_n436_), .A4(new_n427_), .ZN(new_n437_));
  AOI211_X1 g236(.A(new_n391_), .B(new_n405_), .C1(new_n431_), .C2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n431_), .A2(new_n437_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n318_), .A2(KEYINPUT32), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT102), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT103), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n402_), .A2(new_n403_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n391_), .B1(new_n441_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n390_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n380_), .A2(new_n375_), .A3(new_n374_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n368_), .A2(new_n371_), .A3(new_n376_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n388_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n390_), .A2(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n445_), .A2(new_n447_), .B1(new_n454_), .B2(new_n326_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n332_), .A2(new_n438_), .B1(new_n440_), .B2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n278_), .A2(new_n279_), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT30), .Z(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT31), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n457_), .B(KEYINPUT30), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n459_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT83), .B(G15gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT82), .B(G43gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(new_n369_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR3_X1    g272(.A1(new_n465_), .A2(new_n466_), .A3(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n202_), .B1(new_n456_), .B2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n391_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n405_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n440_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n391_), .B1(new_n431_), .B2(new_n437_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n405_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n326_), .A2(KEYINPUT104), .A3(new_n327_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT104), .B1(new_n326_), .B2(new_n327_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n481_), .B(new_n482_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n455_), .A2(new_n440_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n476_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT105), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n477_), .A2(new_n480_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT64), .B(G106gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT10), .B(G99gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G85gat), .B(G92gat), .Z(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(KEYINPUT9), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT6), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT9), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G85gat), .A3(G92gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n497_), .B1(KEYINPUT7), .B2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT65), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n494_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n500_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G29gat), .B(G36gat), .Z(new_n509_));
  XOR2_X1   g308(.A(G43gat), .B(G50gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n505_), .A2(new_n506_), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n508_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n517_));
  NAND2_X1  g316(.A1(G232gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT35), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(KEYINPUT72), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(KEYINPUT35), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n508_), .A2(new_n513_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n511_), .B(KEYINPUT15), .ZN(new_n524_));
  AOI211_X1 g323(.A(new_n521_), .B(new_n522_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n516_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(KEYINPUT72), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(new_n527_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT73), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n516_), .A2(new_n525_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n527_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT73), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT36), .Z(new_n539_));
  NAND3_X1  g338(.A1(new_n531_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n490_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(KEYINPUT106), .Z(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  XOR2_X1   g345(.A(G57gat), .B(G64gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT66), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n549_));
  XOR2_X1   g348(.A(G71gat), .B(G78gat), .Z(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n523_), .A2(new_n546_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n523_), .B(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n556_), .A2(G230gat), .A3(G233gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(G120gat), .B(G148gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n559_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n565_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(KEYINPUT68), .A3(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT13), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n572_), .B1(KEYINPUT69), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT74), .B1(new_n581_), .B2(KEYINPUT17), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G15gat), .B(G22gat), .ZN(new_n583_));
  INV_X1    g382(.A(G1gat), .ZN(new_n584_));
  INV_X1    g383(.A(G8gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT14), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G1gat), .B(G8gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n582_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(new_n554_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n581_), .A2(KEYINPUT17), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n593_), .B2(new_n554_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n524_), .A2(new_n590_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT76), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n589_), .B2(new_n511_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n589_), .A2(new_n511_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT75), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n590_), .A2(new_n512_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n599_), .A2(new_n602_), .B1(new_n606_), .B2(new_n601_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G169gat), .B(G197gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  OR2_X1    g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n610_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n577_), .A2(new_n597_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n545_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n391_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n597_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n476_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n332_), .A2(new_n440_), .A3(new_n482_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n621_), .A2(KEYINPUT105), .B1(new_n623_), .B2(new_n478_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n614_), .B1(new_n624_), .B2(new_n477_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n533_), .A2(new_n539_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n542_), .A2(KEYINPUT37), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n543_), .B2(new_n629_), .ZN(new_n630_));
  AND4_X1   g429(.A1(new_n620_), .A2(new_n625_), .A3(new_n576_), .A4(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n584_), .A3(new_n391_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT38), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n619_), .A2(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n479_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(new_n585_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n616_), .A2(new_n635_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(G8gat), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT39), .B(new_n585_), .C1(new_n616_), .C2(new_n635_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n641_), .B(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n631_), .A2(new_n645_), .A3(new_n476_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G15gat), .B1(new_n617_), .B2(new_n488_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n631_), .A2(new_n652_), .A3(new_n439_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G22gat), .B1(new_n617_), .B2(new_n440_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(G1327gat));
  AND2_X1   g457(.A1(new_n540_), .A2(new_n542_), .ZN(new_n659_));
  AND4_X1   g458(.A1(new_n659_), .A2(new_n625_), .A3(new_n576_), .A4(new_n597_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n391_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n576_), .A2(new_n597_), .A3(new_n613_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n627_), .B1(new_n659_), .B2(KEYINPUT37), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n490_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n490_), .B2(new_n664_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT110), .B(new_n666_), .C1(new_n490_), .C2(new_n664_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT44), .B(new_n662_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT111), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n630_), .B1(new_n624_), .B2(new_n477_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT110), .B1(new_n673_), .B2(new_n666_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n667_), .A2(new_n668_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n665_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(KEYINPUT44), .A4(new_n662_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n662_), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n672_), .A2(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n391_), .A2(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n661_), .B1(new_n681_), .B2(new_n682_), .ZN(G1328gat));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n660_), .A2(new_n684_), .A3(new_n635_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT45), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n672_), .A2(new_n678_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n479_), .B1(new_n680_), .B2(new_n679_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT112), .B1(new_n689_), .B2(G36gat), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT112), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n691_), .B(new_n684_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n686_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI221_X1 g494(.A(new_n686_), .B1(KEYINPUT113), .B2(KEYINPUT46), .C1(new_n690_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  NAND3_X1  g496(.A1(new_n681_), .A2(G43gat), .A3(new_n476_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G43gat), .B1(new_n660_), .B2(new_n476_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT114), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n701_), .B(new_n702_), .Z(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n660_), .B2(new_n439_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n439_), .A2(G50gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n681_), .B2(new_n705_), .ZN(G1331gat));
  INV_X1    g505(.A(G57gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n597_), .A2(new_n613_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n545_), .A2(new_n577_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n709_), .B2(new_n391_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n576_), .A2(new_n597_), .A3(new_n664_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n613_), .B1(new_n624_), .B2(new_n477_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(G57gat), .A3(new_n618_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n710_), .A2(new_n714_), .ZN(G1332gat));
  INV_X1    g514(.A(G64gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n709_), .B2(new_n635_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT48), .Z(new_n718_));
  INV_X1    g517(.A(new_n713_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n716_), .A3(new_n635_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1333gat));
  INV_X1    g520(.A(G71gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n709_), .B2(new_n476_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT49), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n722_), .A3(new_n476_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1334gat));
  INV_X1    g525(.A(G78gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n709_), .B2(new_n439_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT50), .Z(new_n729_));
  NAND3_X1  g528(.A1(new_n719_), .A2(new_n727_), .A3(new_n439_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1335gat));
  AND4_X1   g530(.A1(new_n597_), .A2(new_n676_), .A3(new_n614_), .A4(new_n577_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n618_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n577_), .A2(new_n659_), .A3(new_n597_), .A4(new_n712_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT116), .ZN(new_n736_));
  INV_X1    g535(.A(G85gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n737_), .A3(new_n391_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n734_), .A2(new_n738_), .ZN(G1336gat));
  OAI21_X1  g538(.A(G92gat), .B1(new_n733_), .B2(new_n479_), .ZN(new_n740_));
  INV_X1    g539(.A(G92gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n741_), .A3(new_n635_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1337gat));
  NOR2_X1   g542(.A1(new_n488_), .A2(new_n492_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n736_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G99gat), .B1(new_n733_), .B2(new_n488_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(new_n751_), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  INV_X1    g552(.A(new_n491_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n736_), .A2(new_n439_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n732_), .A2(new_n439_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT53), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n755_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1339gat));
  XNOR2_X1  g563(.A(new_n708_), .B(KEYINPUT118), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n576_), .A2(new_n630_), .A3(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT54), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n599_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n610_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n606_), .A2(new_n600_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT119), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(KEYINPUT119), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n612_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT121), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n566_), .A3(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n612_), .A3(new_n773_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n559_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT121), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n559_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n558_), .B2(new_n557_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n565_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n559_), .B2(new_n781_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n785_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n780_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n630_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n790_), .B2(new_n789_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n613_), .B(new_n566_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n570_), .A2(new_n571_), .A3(new_n774_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n659_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n795_), .A2(KEYINPUT57), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n597_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n767_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n622_), .A2(new_n488_), .A3(new_n618_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT122), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n803_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT120), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n792_), .A3(new_n796_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n795_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n597_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n805_), .B1(new_n809_), .B2(new_n767_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n804_), .B1(new_n810_), .B2(new_n801_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n614_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n810_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n614_), .A2(G113gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(G1340gat));
  OAI21_X1  g614(.A(G120gat), .B1(new_n811_), .B2(new_n576_), .ZN(new_n816_));
  INV_X1    g615(.A(G120gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n576_), .B2(KEYINPUT60), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(KEYINPUT60), .B2(new_n817_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n813_), .B2(new_n819_), .ZN(G1341gat));
  OAI21_X1  g619(.A(G127gat), .B1(new_n811_), .B2(new_n597_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n597_), .A2(G127gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n813_), .B2(new_n822_), .ZN(G1342gat));
  OAI211_X1 g622(.A(new_n804_), .B(new_n664_), .C1(new_n810_), .C2(new_n801_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G134gat), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n813_), .A2(G134gat), .A3(new_n543_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT123), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n826_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n809_), .A2(new_n767_), .ZN(new_n832_));
  NOR4_X1   g631(.A1(new_n635_), .A2(new_n476_), .A3(new_n618_), .A4(new_n440_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n613_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT125), .B1(new_n834_), .B2(new_n614_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT124), .B(G141gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n835_), .A2(new_n577_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g645(.A1(new_n834_), .A2(new_n597_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT61), .B(G155gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  OR3_X1    g648(.A1(new_n834_), .A2(G162gat), .A3(new_n543_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G162gat), .B1(new_n834_), .B2(new_n630_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1347gat));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n439_), .B1(new_n767_), .B2(new_n799_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n488_), .A2(new_n391_), .A3(new_n479_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n614_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n857_), .B2(new_n263_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT62), .B(G169gat), .C1(new_n856_), .C2(new_n614_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(G1348gat));
  INV_X1    g660(.A(new_n856_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G176gat), .B1(new_n862_), .B2(new_n577_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n832_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n439_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n577_), .A2(G176gat), .A3(new_n855_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  AND2_X1   g666(.A1(new_n855_), .A2(new_n620_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G183gat), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n250_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n854_), .B2(new_n871_), .ZN(G1350gat));
  OAI21_X1  g671(.A(G190gat), .B1(new_n856_), .B2(new_n630_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n659_), .A2(new_n252_), .A3(new_n284_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n856_), .B2(new_n874_), .ZN(G1351gat));
  NAND3_X1  g674(.A1(new_n635_), .A2(new_n488_), .A3(new_n481_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n864_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n613_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g678(.A(G204gat), .B1(new_n877_), .B2(new_n577_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n864_), .A2(new_n214_), .A3(new_n576_), .A4(new_n876_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT126), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n877_), .A2(new_n226_), .A3(new_n577_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n864_), .A2(new_n576_), .A3(new_n876_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n883_), .B(new_n884_), .C1(G204gat), .C2(new_n885_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n882_), .A2(new_n886_), .ZN(G1353gat));
  NAND2_X1  g686(.A1(new_n877_), .A2(new_n620_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  AND2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n888_), .B2(new_n889_), .ZN(G1354gat));
  NOR4_X1   g691(.A1(new_n864_), .A2(G218gat), .A3(new_n543_), .A4(new_n876_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT127), .ZN(new_n895_));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n864_), .A2(new_n630_), .A3(new_n876_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n894_), .B(new_n895_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n896_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT127), .B1(new_n899_), .B2(new_n893_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1355gat));
endmodule


