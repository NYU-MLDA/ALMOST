//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G225gat), .A2(G233gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT84), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT3), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(KEYINPUT3), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n217_), .B(KEYINPUT85), .Z(new_n218_));
  OAI211_X1 g017(.A(new_n208_), .B(new_n209_), .C1(new_n216_), .C2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n209_), .B(KEYINPUT1), .Z(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n208_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224_));
  XOR2_X1   g023(.A(G113gat), .B(G120gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n219_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT4), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n223_), .A2(new_n231_), .A3(new_n227_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n206_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n206_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n234_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n205_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT95), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT33), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT95), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(new_n205_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT96), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT33), .B1(new_n236_), .B2(KEYINPUT95), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(KEYINPUT96), .A3(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G226gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT19), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT23), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(G183gat), .B2(G190gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT80), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n250_), .B(new_n254_), .C1(G183gat), .C2(G190gat), .ZN(new_n255_));
  INV_X1    g054(.A(G176gat), .ZN(new_n256_));
  INV_X1    g055(.A(G169gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT22), .B1(new_n257_), .B2(KEYINPUT79), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n257_), .A2(KEYINPUT22), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n256_), .B(new_n258_), .C1(new_n259_), .C2(KEYINPUT79), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .A4(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT25), .B(G183gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n256_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n253_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n265_), .A2(KEYINPUT24), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n250_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G211gat), .B(G218gat), .Z(new_n272_));
  INV_X1    g071(.A(KEYINPUT21), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(KEYINPUT21), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n275_), .B1(new_n276_), .B2(new_n272_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT20), .B1(new_n271_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n267_), .B(KEYINPUT90), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n269_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT22), .B(G169gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n256_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n253_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n251_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n277_), .B1(new_n283_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n248_), .B1(new_n279_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n271_), .A2(new_n278_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n248_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n283_), .A2(new_n289_), .A3(new_n277_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n292_), .B(new_n294_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n295_), .A2(new_n296_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n291_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT18), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G64gat), .B(G92gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n230_), .A2(new_n206_), .A3(new_n232_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n205_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n228_), .A2(new_n229_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n306_), .B(new_n307_), .C1(new_n206_), .C2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n291_), .B(new_n303_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT33), .B(new_n205_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT94), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n312_), .A2(new_n313_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n311_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n246_), .A2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n299_), .A2(new_n319_), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n233_), .A2(new_n205_), .A3(new_n235_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n236_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n295_), .A2(KEYINPUT20), .A3(new_n292_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n248_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n279_), .A2(new_n290_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(new_n248_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n319_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n320_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n318_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT97), .ZN(new_n330_));
  INV_X1    g129(.A(new_n223_), .ZN(new_n331_));
  XOR2_X1   g130(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n332_));
  OAI21_X1  g131(.A(new_n278_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(G228gat), .A3(G233gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n223_), .A2(KEYINPUT29), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT86), .Z(new_n338_));
  NOR2_X1   g137(.A1(new_n277_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n334_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n223_), .A2(KEYINPUT29), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n335_), .A2(new_n339_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT87), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n340_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n346_), .A3(new_n334_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G78gat), .B(G106gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT89), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G22gat), .B(G50gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n348_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n329_), .A2(new_n330_), .A3(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n322_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT98), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n305_), .A2(new_n310_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n326_), .A2(new_n304_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(KEYINPUT27), .A3(new_n310_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n363_), .A2(new_n364_), .A3(new_n367_), .A4(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n369_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n348_), .A2(new_n352_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n356_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n322_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n357_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT98), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n370_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n328_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n246_), .B2(new_n317_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT97), .B1(new_n380_), .B2(new_n360_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n362_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G15gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n271_), .B(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G71gat), .B(G99gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT82), .B(G43gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n385_), .B(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n226_), .B(KEYINPUT31), .Z(new_n392_));
  OR3_X1    g191(.A1(new_n391_), .A2(KEYINPUT83), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(KEYINPUT83), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n392_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n391_), .A2(KEYINPUT83), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n371_), .A2(KEYINPUT99), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT99), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n367_), .A2(new_n399_), .A3(new_n369_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n397_), .A2(new_n322_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n361_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT100), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n401_), .A2(KEYINPUT100), .A3(new_n361_), .A4(new_n402_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n382_), .A2(new_n397_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G1gat), .B(G8gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT77), .ZN(new_n409_));
  INV_X1    g208(.A(G15gat), .ZN(new_n410_));
  INV_X1    g209(.A(G22gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G15gat), .A2(G22gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G1gat), .A2(G8gat), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n412_), .A2(new_n413_), .B1(KEYINPUT14), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n409_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G29gat), .B(G36gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(KEYINPUT74), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(G36gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G29gat), .ZN(new_n421_));
  INV_X1    g220(.A(G29gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G36gat), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n421_), .A2(new_n423_), .A3(KEYINPUT74), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G43gat), .B(G50gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n416_), .B(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(G229gat), .A3(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n416_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n430_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G229gat), .A2(G233gat), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n427_), .A2(new_n429_), .A3(KEYINPUT15), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT15), .B1(new_n427_), .B2(new_n429_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n435_), .B(new_n436_), .C1(new_n440_), .C2(new_n434_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n433_), .A2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G113gat), .B(G141gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT78), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G169gat), .B(G197gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n433_), .A2(new_n441_), .A3(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G230gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G78gat), .ZN(new_n456_));
  INV_X1    g255(.A(G78gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n457_), .A3(new_n454_), .ZN(new_n458_));
  INV_X1    g257(.A(G64gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G57gat), .ZN(new_n460_));
  INV_X1    g259(.A(G57gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G64gat), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n460_), .A2(new_n462_), .A3(KEYINPUT11), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT11), .B1(new_n460_), .B2(new_n462_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n456_), .B(new_n458_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n460_), .A2(new_n462_), .A3(KEYINPUT11), .ZN(new_n466_));
  INV_X1    g265(.A(new_n458_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n457_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT9), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(KEYINPUT6), .ZN(new_n484_));
  OAI22_X1  g283(.A1(new_n482_), .A2(new_n484_), .B1(KEYINPUT9), .B2(new_n478_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT64), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n478_), .A2(KEYINPUT9), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(KEYINPUT6), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n474_), .A4(new_n479_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  AND2_X1   g293(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n488_), .A2(new_n489_), .ZN(new_n498_));
  OR2_X1    g297(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n499_));
  INV_X1    g298(.A(G99gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n472_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n477_), .A2(new_n478_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n493_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(KEYINPUT8), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT66), .B1(new_n482_), .B2(new_n484_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n488_), .A2(new_n489_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT67), .B1(new_n497_), .B2(new_n502_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n497_), .A2(new_n502_), .A3(KEYINPUT67), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n509_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n470_), .B1(new_n508_), .B2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n518_), .A2(KEYINPUT69), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n486_), .A2(new_n492_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n488_), .A2(new_n489_), .A3(new_n511_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n511_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n501_), .B1(new_n525_), .B2(new_n499_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n494_), .A2(new_n496_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n524_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n523_), .A2(new_n528_), .A3(new_n516_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n509_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n470_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n520_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n518_), .B2(KEYINPUT69), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n452_), .B1(new_n519_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n518_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n520_), .A2(new_n531_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n470_), .A2(KEYINPUT70), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n465_), .A2(new_n469_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n542_), .A3(KEYINPUT12), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n537_), .A2(new_n451_), .A3(new_n543_), .A4(new_n533_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n535_), .A2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G120gat), .B(G148gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT5), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n545_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT71), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n550_), .B2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n556_), .A2(KEYINPUT72), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(KEYINPUT72), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n450_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n407_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT75), .B1(new_n439_), .B2(new_n538_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT73), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n439_), .B2(new_n538_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n520_), .A2(new_n531_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n430_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n572_), .B(new_n574_), .C1(new_n565_), .C2(new_n569_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n564_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n578_), .A3(new_n577_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT76), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n581_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n416_), .B(new_n592_), .Z(new_n593_));
  AOI211_X1 g392(.A(new_n587_), .B(new_n591_), .C1(new_n593_), .C2(new_n542_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n593_), .B2(new_n542_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n591_), .B(new_n587_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n593_), .B2(new_n532_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n593_), .B2(new_n532_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n586_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n560_), .A2(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n601_), .A2(G1gat), .A3(new_n375_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT102), .Z(new_n605_));
  NOR2_X1   g404(.A1(new_n602_), .A2(new_n603_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT103), .ZN(new_n607_));
  INV_X1    g406(.A(new_n599_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n581_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n407_), .A2(new_n559_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n375_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n605_), .A2(new_n607_), .A3(new_n613_), .ZN(G1324gat));
  NAND2_X1  g413(.A1(new_n382_), .A2(new_n397_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n405_), .A2(new_n406_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n559_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n401_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n610_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .A4(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n621_), .A2(new_n622_), .A3(G8gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n621_), .B2(G8gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT39), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(G8gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT104), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n621_), .A2(new_n622_), .A3(G8gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT105), .B(KEYINPUT39), .C1(new_n623_), .C2(new_n624_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n629_), .A2(KEYINPUT106), .A3(new_n630_), .A4(new_n631_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n627_), .A2(new_n634_), .A3(new_n635_), .A4(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n601_), .ZN(new_n638_));
  INV_X1    g437(.A(G8gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n619_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n637_), .A2(KEYINPUT40), .A3(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  INV_X1    g444(.A(new_n397_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n410_), .B1(new_n611_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n638_), .A2(new_n410_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  AOI21_X1  g450(.A(new_n411_), .B1(new_n611_), .B2(new_n360_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n638_), .A2(new_n411_), .A3(new_n360_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  NOR2_X1   g455(.A1(new_n608_), .A2(new_n609_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n560_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n322_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n617_), .A2(new_n660_), .A3(new_n586_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n586_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n407_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n599_), .A3(new_n618_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n664_), .A2(KEYINPUT44), .A3(new_n599_), .A4(new_n618_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n375_), .A2(new_n422_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n659_), .B1(new_n669_), .B2(new_n670_), .ZN(G1328gat));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n668_), .A3(new_n619_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G36gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n658_), .A2(new_n420_), .A3(new_n619_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1329gat));
  NAND3_X1  g477(.A1(new_n669_), .A2(G43gat), .A3(new_n646_), .ZN(new_n679_));
  INV_X1    g478(.A(G43gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n658_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n397_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(new_n685_), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  OR3_X1    g486(.A1(new_n681_), .A2(G50gat), .A3(new_n361_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n669_), .A2(new_n689_), .A3(new_n360_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n669_), .B2(new_n360_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(G1331gat));
  NOR2_X1   g492(.A1(new_n557_), .A2(new_n558_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n450_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n407_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n600_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n461_), .A3(new_n322_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n697_), .A2(new_n407_), .A3(new_n610_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n322_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n461_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT110), .ZN(G1332gat));
  AOI21_X1  g503(.A(new_n459_), .B1(new_n701_), .B2(new_n619_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT48), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n699_), .A2(new_n459_), .A3(new_n619_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n701_), .B2(new_n646_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT49), .Z(new_n711_));
  NAND2_X1  g510(.A1(new_n646_), .A2(new_n709_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT111), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n699_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1334gat));
  AOI21_X1  g514(.A(new_n457_), .B1(new_n701_), .B2(new_n360_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n457_), .A3(new_n360_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1335gat));
  NAND3_X1  g519(.A1(new_n664_), .A2(new_n599_), .A3(new_n696_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721_), .B2(new_n375_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n698_), .A2(new_n657_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n475_), .A3(new_n322_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1336gat));
  OAI21_X1  g525(.A(G92gat), .B1(new_n721_), .B2(new_n401_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(new_n476_), .A3(new_n619_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1337gat));
  OAI21_X1  g528(.A(G99gat), .B1(new_n721_), .B2(new_n397_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n724_), .A2(new_n471_), .A3(new_n473_), .A4(new_n646_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT113), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n472_), .A3(new_n360_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n664_), .A2(new_n599_), .A3(new_n360_), .A4(new_n696_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G106gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G106gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1339gat));
  NAND2_X1  g540(.A1(new_n450_), .A2(G113gat), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT119), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n450_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n600_), .A2(new_n745_), .A3(new_n556_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT54), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n545_), .A2(new_n549_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n450_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT115), .B1(new_n544_), .B2(new_n750_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n465_), .A2(new_n469_), .A3(new_n540_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n540_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT12), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n533_), .B1(new_n573_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT12), .B1(new_n538_), .B2(new_n470_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(KEYINPUT55), .A4(new_n451_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n751_), .A2(new_n759_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n755_), .A2(new_n452_), .A3(new_n756_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n537_), .A2(new_n543_), .A3(new_n533_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n452_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n763_), .B2(KEYINPUT55), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n549_), .B1(new_n760_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n750_), .B1(new_n762_), .B2(new_n452_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n751_), .B(new_n759_), .C1(new_n768_), .C2(new_n761_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n549_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n749_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n446_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n435_), .B1(new_n440_), .B2(new_n434_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n436_), .B2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(new_n449_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n550_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT57), .B(new_n609_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n748_), .A2(new_n775_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n586_), .B1(new_n780_), .B2(KEYINPUT58), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n782_), .B(new_n779_), .C1(new_n767_), .C2(new_n770_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n749_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n770_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n549_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n581_), .B1(new_n788_), .B2(new_n776_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(KEYINPUT57), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n599_), .B1(new_n784_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n747_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NOR4_X1   g592(.A1(new_n619_), .A2(new_n397_), .A3(new_n375_), .A4(new_n360_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n789_), .B2(KEYINPUT57), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n771_), .A2(new_n777_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT116), .B(new_n798_), .C1(new_n799_), .C2(new_n581_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n784_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n599_), .B1(new_n801_), .B2(KEYINPUT117), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n784_), .C1(new_n797_), .C2(new_n800_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n747_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT118), .B(new_n747_), .C1(new_n802_), .C2(new_n804_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n794_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n744_), .B(new_n795_), .C1(new_n809_), .C2(KEYINPUT59), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n807_), .A2(new_n450_), .A3(new_n808_), .A4(new_n794_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT120), .B1(new_n810_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n795_), .B1(new_n809_), .B2(KEYINPUT59), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n743_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n813_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(new_n809_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT60), .ZN(new_n822_));
  AOI21_X1  g621(.A(G120gat), .B1(new_n694_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT121), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n822_), .B2(G120gat), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n821_), .B(new_n824_), .C1(new_n823_), .C2(new_n826_), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n695_), .B(new_n795_), .C1(new_n809_), .C2(KEYINPUT59), .ZN(new_n828_));
  OAI21_X1  g627(.A(G120gat), .B1(new_n828_), .B2(KEYINPUT122), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n816_), .A2(KEYINPUT122), .A3(new_n694_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(G1341gat));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n821_), .A2(new_n832_), .A3(new_n608_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n816_), .A2(new_n608_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n832_), .ZN(G1342gat));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836_));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n816_), .B2(new_n586_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n809_), .A2(G134gat), .A3(new_n609_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n836_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n662_), .B(new_n795_), .C1(new_n809_), .C2(KEYINPUT59), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(KEYINPUT123), .C1(new_n842_), .C2(new_n837_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(G1343gat));
  AND2_X1   g643(.A1(new_n807_), .A2(new_n808_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n397_), .A2(new_n360_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n619_), .A2(new_n375_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n745_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT124), .B(G141gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n848_), .A2(new_n695_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT125), .B(G148gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NOR2_X1   g653(.A1(new_n848_), .A2(new_n599_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT61), .B(G155gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  OAI21_X1  g656(.A(G162gat), .B1(new_n848_), .B2(new_n662_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n609_), .A2(G162gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n848_), .B2(new_n859_), .ZN(G1347gat));
  NAND2_X1  g659(.A1(new_n619_), .A2(new_n402_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n360_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n792_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n257_), .B1(new_n864_), .B2(new_n450_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n865_), .A2(KEYINPUT62), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(KEYINPUT62), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n450_), .A3(new_n284_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT126), .ZN(G1348gat));
  AOI21_X1  g669(.A(G176gat), .B1(new_n864_), .B2(new_n694_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n845_), .A2(new_n361_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n695_), .A2(new_n256_), .A3(new_n861_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  NOR3_X1   g673(.A1(new_n863_), .A2(new_n599_), .A3(new_n262_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT127), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n872_), .A2(new_n608_), .A3(new_n619_), .A4(new_n402_), .ZN(new_n877_));
  INV_X1    g676(.A(G183gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n863_), .B2(new_n662_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n581_), .A2(new_n263_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n863_), .B2(new_n881_), .ZN(G1351gat));
  NOR3_X1   g681(.A1(new_n401_), .A2(new_n846_), .A3(new_n322_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n845_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n450_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n694_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g687(.A1(new_n845_), .A2(new_n608_), .A3(new_n883_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  AND2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n889_), .B2(new_n890_), .ZN(G1354gat));
  INV_X1    g692(.A(new_n884_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G218gat), .B1(new_n894_), .B2(new_n662_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n609_), .A2(G218gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(new_n896_), .ZN(G1355gat));
endmodule


