//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n208_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G229gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n216_));
  XNOR2_X1  g015(.A(new_n211_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n208_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(new_n211_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n213_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G141gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G169gat), .B(G197gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n223_), .B(new_n224_), .Z(new_n225_));
  XOR2_X1   g024(.A(new_n222_), .B(new_n225_), .Z(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT76), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT22), .ZN(new_n231_));
  AOI21_X1  g030(.A(G176gat), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n228_), .B(KEYINPUT22), .C1(new_n230_), .C2(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(KEYINPUT78), .A3(new_n235_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240_));
  INV_X1    g039(.A(G183gat), .ZN(new_n241_));
  INV_X1    g040(.A(G190gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n243_), .B(new_n244_), .C1(G183gat), .C2(G190gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n238_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n244_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(KEYINPUT24), .A3(new_n235_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT75), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT25), .B(G183gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n242_), .A2(KEYINPUT26), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(KEYINPUT75), .B2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n250_), .B(new_n252_), .C1(new_n255_), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n246_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT80), .ZN(new_n263_));
  XOR2_X1   g062(.A(G127gat), .B(G134gat), .Z(new_n264_));
  INV_X1    g063(.A(G120gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G113gat), .ZN(new_n266_));
  INV_X1    g065(.A(G113gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G120gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n272_), .A3(KEYINPUT82), .ZN(new_n273_));
  OR3_X1    g072(.A1(new_n264_), .A2(new_n269_), .A3(KEYINPUT82), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n275_), .A2(KEYINPUT31), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(KEYINPUT31), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT81), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n263_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n262_), .A2(KEYINPUT80), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281_));
  INV_X1    g080(.A(G43gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G15gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n279_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n290_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(KEYINPUT21), .ZN(new_n297_));
  INV_X1    g096(.A(G197gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT21), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(new_n290_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n295_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT90), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G228gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT86), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(KEYINPUT85), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n311_), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n307_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT87), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT2), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G141gat), .A3(G148gat), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n315_), .A2(new_n317_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n309_), .A2(KEYINPUT85), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n311_), .B1(G141gat), .B2(G148gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n323_), .A2(KEYINPUT86), .A3(new_n324_), .A4(new_n308_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n313_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n326_));
  OR3_X1    g125(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n327_), .A2(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n333_), .A3(new_n331_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT1), .B1(new_n335_), .B2(new_n329_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n328_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n309_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n339_), .A2(new_n318_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n326_), .A2(new_n332_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n304_), .B(new_n305_), .C1(new_n306_), .C2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n306_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n294_), .B1(new_n291_), .B2(new_n290_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT21), .B(new_n299_), .C1(new_n296_), .C2(KEYINPUT89), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n344_), .A2(new_n345_), .B1(new_n294_), .B2(new_n292_), .ZN(new_n346_));
  OAI211_X1 g145(.A(G228gat), .B(G233gat), .C1(new_n343_), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G78gat), .B(G106gat), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(new_n347_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n326_), .A2(new_n332_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n338_), .A2(new_n340_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G22gat), .B(G50gat), .Z(new_n357_));
  NOR3_X1   g156(.A1(new_n356_), .A2(KEYINPUT29), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n359_));
  INV_X1    g158(.A(new_n357_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n341_), .B2(new_n306_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n353_), .A2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n350_), .A2(new_n362_), .A3(new_n363_), .A4(new_n352_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT100), .ZN(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT98), .ZN(new_n370_));
  XOR2_X1   g169(.A(G1gat), .B(G29gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G57gat), .B(G85gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n273_), .A2(new_n274_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n356_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT95), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n356_), .A2(new_n381_), .A3(new_n376_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT95), .B1(new_n341_), .B2(new_n275_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n270_), .A2(new_n272_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n354_), .A2(new_n355_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n382_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT4), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT96), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(KEYINPUT96), .A3(KEYINPUT4), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n380_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n378_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n374_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n380_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n354_), .A2(new_n355_), .A3(new_n384_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n396_), .B(KEYINPUT95), .C1(new_n341_), .C2(new_n275_), .ZN(new_n397_));
  AOI211_X1 g196(.A(new_n388_), .B(new_n375_), .C1(new_n397_), .C2(new_n382_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT96), .B1(new_n386_), .B2(KEYINPUT4), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n395_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n393_), .A2(new_n374_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n400_), .A2(KEYINPUT99), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT99), .B1(new_n400_), .B2(new_n401_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n394_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT22), .B(G169gat), .ZN(new_n406_));
  INV_X1    g205(.A(G176gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n245_), .A2(new_n235_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n235_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT93), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT93), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n413_), .A3(new_n235_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n251_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n410_), .A2(new_n251_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n247_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n253_), .A2(new_n256_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n409_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n405_), .B1(new_n421_), .B2(new_n303_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n304_), .B2(new_n260_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT19), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT91), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n304_), .A2(new_n260_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n409_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n420_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(new_n415_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n405_), .B1(new_n432_), .B2(new_n346_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G8gat), .B(G36gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n427_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n423_), .A2(new_n426_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n429_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n445_), .B2(new_n441_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n368_), .B1(new_n404_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n434_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n426_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n346_), .A2(KEYINPUT90), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n303_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n259_), .A3(new_n246_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n455_), .B2(new_n422_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n439_), .B1(new_n449_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n427_), .A2(new_n434_), .A3(new_n440_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n378_), .B(new_n377_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n374_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n386_), .B2(new_n379_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n400_), .A2(KEYINPUT33), .A3(new_n401_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n392_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n391_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n463_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n448_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n404_), .A2(new_n368_), .A3(new_n447_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n367_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n367_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT27), .B1(new_n457_), .B2(new_n458_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n439_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n474_), .A2(KEYINPUT27), .A3(new_n458_), .ZN(new_n475_));
  NOR4_X1   g274(.A1(new_n404_), .A2(new_n472_), .A3(new_n473_), .A4(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n289_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n461_), .B1(new_n400_), .B2(new_n392_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT99), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n391_), .B2(new_n466_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n400_), .A2(KEYINPUT99), .A3(new_n401_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n478_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n288_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT102), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT101), .B1(new_n475_), .B2(new_n473_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT27), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n459_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT101), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n474_), .A2(KEYINPUT27), .A3(new_n458_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n485_), .B1(new_n492_), .B2(new_n472_), .ZN(new_n493_));
  AOI211_X1 g292(.A(KEYINPUT102), .B(new_n367_), .C1(new_n486_), .C2(new_n491_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n484_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n227_), .B1(new_n477_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT10), .B(G99gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(G106gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT65), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT6), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(G99gat), .A3(G106gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT66), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n505_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G85gat), .ZN(new_n512_));
  INV_X1    g311(.A(G92gat), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT9), .ZN(new_n514_));
  XOR2_X1   g313(.A(G85gat), .B(G92gat), .Z(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(KEYINPUT9), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n501_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n515_), .B1(new_n520_), .B2(new_n506_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT8), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n515_), .A2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G71gat), .B(G78gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n528_), .B1(KEYINPUT11), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n529_), .A2(new_n531_), .A3(KEYINPUT11), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n529_), .B2(KEYINPUT11), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n530_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n527_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n517_), .A3(new_n526_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(KEYINPUT12), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n527_), .A2(new_n537_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(KEYINPUT64), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n538_), .A2(new_n539_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n545_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n545_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n554_), .B(KEYINPUT69), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT13), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(KEYINPUT13), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT70), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT74), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n208_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(new_n536_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n536_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n569_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n517_), .A2(new_n526_), .A3(new_n211_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT72), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT34), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n527_), .A2(new_n217_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n581_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT73), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n586_), .A2(new_n590_), .A3(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n580_), .A2(new_n591_), .A3(new_n587_), .A4(new_n585_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT36), .Z(new_n599_));
  AND3_X1   g398(.A1(new_n594_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(KEYINPUT36), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT37), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  AOI211_X1 g403(.A(new_n589_), .B(new_n592_), .C1(new_n580_), .C2(new_n585_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n595_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n601_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n594_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n577_), .A2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n497_), .A2(new_n564_), .A3(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n203_), .A3(new_n404_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n600_), .A2(new_n603_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n477_), .B2(new_n495_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n562_), .A2(new_n226_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n577_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n482_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n614_), .A2(new_n615_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n616_), .A2(new_n623_), .A3(new_n624_), .ZN(G1324gat));
  OAI21_X1  g424(.A(G8gat), .B1(new_n622_), .B2(new_n492_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT39), .ZN(new_n627_));
  INV_X1    g426(.A(new_n492_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n613_), .A2(new_n204_), .A3(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n622_), .B2(new_n289_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  INV_X1    g432(.A(new_n613_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(G15gat), .A3(new_n289_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1326gat));
  OAI21_X1  g435(.A(G22gat), .B1(new_n622_), .B2(new_n472_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT42), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n472_), .A2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n634_), .B2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n619_), .A2(new_n577_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT100), .B1(new_n482_), .B2(new_n446_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n463_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n470_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n476_), .B1(new_n644_), .B2(new_n472_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n495_), .B1(new_n645_), .B2(new_n288_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n611_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT43), .B1(new_n611_), .B2(KEYINPUT103), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n641_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT44), .B(new_n641_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n404_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G29gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n620_), .A2(new_n617_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n562_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n496_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n482_), .A2(G29gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n661_), .B2(new_n662_), .ZN(G1328gat));
  NOR2_X1   g462(.A1(new_n492_), .A2(G36gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n496_), .A2(new_n659_), .A3(new_n664_), .A4(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n646_), .A2(new_n226_), .A3(new_n659_), .A4(new_n664_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n666_), .A2(new_n667_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n667_), .B1(new_n666_), .B2(new_n670_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(KEYINPUT107), .A2(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n653_), .A2(new_n628_), .A3(new_n654_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(KEYINPUT104), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n653_), .A2(new_n678_), .A3(new_n628_), .A4(new_n654_), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT46), .B(new_n674_), .C1(new_n677_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(KEYINPUT104), .ZN(new_n682_));
  INV_X1    g481(.A(new_n675_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n679_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n674_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n680_), .A2(new_n686_), .ZN(G1329gat));
  NAND4_X1  g486(.A1(new_n653_), .A2(G43gat), .A3(new_n288_), .A4(new_n654_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n282_), .B1(new_n661_), .B2(new_n289_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g490(.A1(new_n661_), .A2(G50gat), .A3(new_n472_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n653_), .A2(new_n367_), .A3(new_n654_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(G50gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n693_), .B2(G50gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(G1331gat));
  AOI21_X1  g496(.A(new_n226_), .B1(new_n477_), .B2(new_n495_), .ZN(new_n698_));
  AND4_X1   g497(.A1(new_n658_), .A2(new_n698_), .A3(new_n577_), .A4(new_n611_), .ZN(new_n699_));
  INV_X1    g498(.A(G57gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n404_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n618_), .A2(new_n227_), .A3(new_n564_), .A4(new_n577_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n482_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1332gat));
  OAI21_X1  g503(.A(G64gat), .B1(new_n702_), .B2(new_n492_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT48), .ZN(new_n706_));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n699_), .A2(new_n707_), .A3(new_n628_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n702_), .B2(new_n289_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT49), .ZN(new_n711_));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n699_), .A2(new_n712_), .A3(new_n288_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1334gat));
  OAI21_X1  g513(.A(G78gat), .B1(new_n702_), .B2(new_n472_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT50), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n472_), .A2(G78gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT109), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n699_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1335gat));
  NAND3_X1  g519(.A1(new_n658_), .A2(new_n620_), .A3(new_n227_), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n649_), .A2(new_n650_), .A3(KEYINPUT110), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT110), .B1(new_n649_), .B2(new_n650_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(new_n404_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n563_), .A2(new_n657_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n698_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n404_), .A2(new_n512_), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n725_), .A2(new_n512_), .B1(new_n727_), .B2(new_n728_), .ZN(G1336gat));
  AND3_X1   g528(.A1(new_n724_), .A2(G92gat), .A3(new_n628_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n513_), .B1(new_n727_), .B2(new_n492_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT111), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n730_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1337gat));
  NOR3_X1   g535(.A1(new_n727_), .A2(new_n289_), .A3(new_n498_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n724_), .A2(new_n288_), .ZN(new_n739_));
  INV_X1    g538(.A(G99gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT51), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n738_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1338gat));
  NOR3_X1   g544(.A1(new_n727_), .A2(G106gat), .A3(new_n472_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n721_), .A2(new_n472_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(G106gat), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT52), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT52), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n493_), .A2(new_n494_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n289_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n617_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n222_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n219_), .A2(new_n220_), .A3(new_n214_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n225_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n760_), .A2(new_n225_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n559_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n226_), .A2(new_n555_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n540_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n547_), .A2(KEYINPUT55), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n558_), .B1(new_n556_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n769_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n765_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n764_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n769_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n769_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n226_), .B(new_n555_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n759_), .B1(new_n776_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n555_), .A2(new_n763_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(KEYINPUT58), .C1(new_n777_), .C2(new_n778_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT116), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n611_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n781_), .A2(new_n782_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n779_), .A2(KEYINPUT114), .B1(new_n559_), .B2(new_n763_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n774_), .A2(new_n775_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n617_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT57), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n577_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n795_));
  AND4_X1   g594(.A1(new_n227_), .A2(new_n562_), .A3(new_n577_), .A4(new_n611_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT54), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n404_), .B(new_n758_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n756_), .B1(new_n798_), .B2(KEYINPUT59), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n756_), .A3(KEYINPUT59), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n798_), .B2(KEYINPUT59), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n785_), .A2(KEYINPUT116), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n785_), .A2(KEYINPUT116), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n789_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n793_), .B2(KEYINPUT57), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n781_), .A2(new_n782_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n620_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n796_), .B(KEYINPUT54), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n482_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n812_), .A2(KEYINPUT118), .A3(new_n813_), .A4(new_n758_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n804_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n802_), .A2(new_n226_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G113gat), .ZN(new_n817_));
  INV_X1    g616(.A(new_n798_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n267_), .A3(new_n226_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(new_n801_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n815_), .B(new_n564_), .C1(new_n799_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n802_), .A2(KEYINPUT119), .A3(new_n564_), .A4(new_n815_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(G120gat), .A3(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n265_), .B1(new_n562_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n818_), .B(new_n827_), .C1(KEYINPUT60), .C2(new_n265_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1341gat));
  AOI21_X1  g628(.A(G127gat), .B1(new_n818_), .B2(new_n577_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n802_), .A2(new_n815_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n577_), .A2(G127gat), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT120), .Z(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(new_n831_), .B2(new_n833_), .ZN(G1342gat));
  NAND3_X1  g633(.A1(new_n802_), .A2(new_n647_), .A3(new_n815_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G134gat), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n759_), .A2(G134gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n798_), .B2(new_n837_), .ZN(G1343gat));
  NOR2_X1   g637(.A1(new_n288_), .A2(new_n472_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n812_), .A2(new_n492_), .A3(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n227_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n563_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT121), .B(G148gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1345gat));
  NOR2_X1   g644(.A1(new_n840_), .A2(new_n620_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT61), .B(G155gat), .Z(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  OAI21_X1  g647(.A(G162gat), .B1(new_n840_), .B2(new_n611_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n759_), .A2(G162gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n840_), .B2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT122), .ZN(G1347gat));
  AOI21_X1  g651(.A(new_n367_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n483_), .A2(new_n492_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n226_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT123), .Z(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G169gat), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n858_), .A2(KEYINPUT62), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(KEYINPUT62), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n853_), .A2(new_n854_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n226_), .A2(new_n406_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n859_), .A2(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI221_X1 g664(.A(KEYINPUT124), .B1(new_n861_), .B2(new_n862_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1348gat));
  OAI21_X1  g666(.A(G176gat), .B1(new_n861_), .B2(new_n563_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n658_), .A2(new_n407_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n861_), .B2(new_n869_), .ZN(G1349gat));
  NOR2_X1   g669(.A1(new_n861_), .A2(new_n620_), .ZN(new_n871_));
  MUX2_X1   g670(.A(G183gat), .B(new_n256_), .S(new_n871_), .Z(G1350gat));
  NAND3_X1  g671(.A1(new_n853_), .A2(new_n647_), .A3(new_n854_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT125), .B1(new_n873_), .B2(G190gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n617_), .A2(new_n253_), .ZN(new_n877_));
  OAI22_X1  g676(.A1(new_n875_), .A2(new_n876_), .B1(new_n861_), .B2(new_n877_), .ZN(G1351gat));
  NAND3_X1  g677(.A1(new_n628_), .A2(new_n839_), .A3(new_n482_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n226_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n564_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT126), .B(G204gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1353gat));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n577_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  AND2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n886_), .B2(new_n887_), .ZN(G1354gat));
  INV_X1    g689(.A(G218gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n880_), .A2(new_n891_), .A3(new_n617_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n880_), .A2(new_n647_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1355gat));
endmodule


