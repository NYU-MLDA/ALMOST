//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT81), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT81), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n211_), .B(new_n216_), .C1(new_n222_), .C2(KEYINPUT24), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT24), .B1(new_n219_), .B2(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n214_), .A2(new_n215_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT82), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(G183gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT25), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT26), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT80), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(G190gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n232_), .A2(KEYINPUT26), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n231_), .B(new_n234_), .C1(new_n238_), .C2(KEYINPUT80), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(G169gat), .B2(G176gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n222_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n223_), .A2(new_n226_), .A3(new_n239_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n229_), .A2(new_n232_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n216_), .A2(KEYINPUT84), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n214_), .A2(new_n244_), .A3(new_n215_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT22), .B1(new_n217_), .B2(KEYINPUT83), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n217_), .A2(KEYINPUT22), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n218_), .B(new_n250_), .C1(new_n251_), .C2(KEYINPUT83), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n245_), .A2(new_n248_), .A3(new_n249_), .A4(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G218gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G211gat), .ZN(new_n255_));
  INV_X1    g054(.A(G211gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G218gat), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n255_), .A2(new_n257_), .A3(KEYINPUT91), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT91), .B1(new_n255_), .B2(new_n257_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n261_));
  INV_X1    g060(.A(G204gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G197gat), .A2(G204gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n261_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n264_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(G204gat), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(KEYINPUT92), .A3(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n260_), .A2(new_n267_), .A3(KEYINPUT21), .A4(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n255_), .A2(new_n257_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT91), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n255_), .A2(new_n257_), .A3(KEYINPUT91), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n263_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n274_), .B1(G197gat), .B2(G204gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n275_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n243_), .A2(new_n253_), .B1(new_n273_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT94), .B1(new_n228_), .B2(new_n230_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT95), .B1(new_n236_), .B2(new_n237_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n229_), .A2(KEYINPUT25), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n227_), .A2(G183gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT94), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n235_), .A2(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n233_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n286_), .A2(new_n287_), .A3(new_n291_), .A4(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n240_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n222_), .B2(new_n241_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT22), .B(G169gat), .Z(new_n300_));
  OAI211_X1 g099(.A(new_n246_), .B(new_n249_), .C1(new_n300_), .C2(G176gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n273_), .A2(new_n299_), .A3(new_n284_), .A4(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT20), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT100), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n285_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n210_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n273_), .A2(new_n284_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n299_), .A2(new_n301_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n243_), .A2(new_n253_), .A3(new_n284_), .A4(new_n273_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT20), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(new_n209_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n207_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT103), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(KEYINPUT103), .B(new_n207_), .C1(new_n307_), .C2(new_n313_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n303_), .A2(new_n285_), .A3(new_n209_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n210_), .B1(new_n320_), .B2(new_n311_), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n318_), .A2(new_n321_), .A3(new_n207_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n312_), .A2(new_n209_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n243_), .A2(new_n253_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n308_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n328_), .A2(KEYINPUT20), .A3(new_n210_), .A4(new_n302_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n206_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n323_), .B1(new_n322_), .B2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(G71gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G99gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n327_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G134gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G127gat), .ZN(new_n341_));
  INV_X1    g140(.A(G127gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G134gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n339_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n341_), .A2(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT86), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n345_), .A3(new_n338_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n337_), .B(new_n352_), .Z(new_n353_));
  XNOR2_X1  g152(.A(G15gat), .B(G43gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT85), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT30), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT31), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n353_), .B(new_n357_), .Z(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G141gat), .B(G148gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(KEYINPUT1), .B2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n364_), .A2(KEYINPUT1), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G141gat), .ZN(new_n368_));
  INV_X1    g167(.A(G148gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(KEYINPUT3), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(G141gat), .B2(G148gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n370_), .A2(new_n372_), .B1(new_n373_), .B2(KEYINPUT87), .ZN(new_n374_));
  AND3_X1   g173(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G155gat), .B(G162gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n367_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n361_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n374_), .B2(new_n380_), .ZN(new_n387_));
  NOR4_X1   g186(.A1(new_n387_), .A2(new_n367_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n360_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n370_), .A2(new_n372_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n373_), .A2(KEYINPUT87), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n373_), .B2(KEYINPUT87), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n383_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n365_), .A2(new_n366_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n362_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n385_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT28), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n384_), .A2(new_n361_), .A3(new_n385_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n359_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n389_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT93), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n389_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT89), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT29), .B1(new_n387_), .B2(new_n367_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n308_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT88), .B(G233gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G228gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n308_), .A2(new_n407_), .A3(new_n408_), .A4(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n404_), .A2(new_n406_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n406_), .B2(new_n417_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n346_), .A2(new_n339_), .A3(new_n347_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n338_), .B1(new_n350_), .B2(new_n345_), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n420_), .A2(new_n421_), .B1(new_n387_), .B2(new_n367_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n395_), .A2(new_n351_), .A3(new_n348_), .A4(new_n398_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT4), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n395_), .A2(new_n398_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n352_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n425_), .B1(new_n426_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G57gat), .B(G85gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G1gat), .B(G29gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G57gat), .B(G85gat), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n440_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n434_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n433_), .A3(new_n443_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n432_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT101), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n446_), .A2(new_n448_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n452_), .B(new_n425_), .C1(new_n426_), .C2(new_n431_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n432_), .A2(KEYINPUT101), .A3(new_n449_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n454_), .A2(KEYINPUT102), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT102), .B1(new_n454_), .B2(new_n455_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n332_), .A2(new_n358_), .A3(new_n419_), .A4(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n417_), .A2(new_n406_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n417_), .A2(new_n406_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n404_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n331_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n458_), .A2(new_n325_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n326_), .A2(new_n465_), .A3(new_n329_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(new_n455_), .A3(new_n454_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n453_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n429_), .A2(new_n424_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n426_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n422_), .A2(new_n423_), .A3(new_n430_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n449_), .A2(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n453_), .A2(new_n470_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n326_), .A2(new_n206_), .A3(new_n329_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n207_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n471_), .A2(new_n476_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n469_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n419_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n358_), .B1(new_n464_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n459_), .B1(new_n482_), .B2(KEYINPUT104), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n462_), .B1(new_n469_), .B2(new_n479_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n331_), .A2(new_n462_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n485_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n484_), .B1(new_n486_), .B2(new_n325_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT104), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n358_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n483_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT9), .ZN(new_n491_));
  INV_X1    g290(.A(G85gat), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n491_), .B(new_n494_), .C1(new_n496_), .C2(KEYINPUT64), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT6), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(KEYINPUT10), .B(G99gat), .Z(new_n503_));
  INV_X1    g302(.A(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n494_), .A2(new_n506_), .A3(KEYINPUT9), .A4(new_n495_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n497_), .A2(new_n502_), .A3(new_n505_), .A4(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510_));
  INV_X1    g309(.A(G99gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n504_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n509_), .B(new_n512_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  INV_X1    g313(.A(new_n496_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n508_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G71gat), .B(G78gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(KEYINPUT11), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n522_));
  INV_X1    g321(.A(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT66), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n517_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n508_), .A4(new_n526_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n526_), .B(new_n508_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT65), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n529_), .A2(new_n531_), .A3(new_n536_), .A4(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(G230gat), .A3(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n528_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n518_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT67), .B(new_n508_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(KEYINPUT12), .A3(new_n547_), .A4(new_n527_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n543_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n540_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G120gat), .B(G148gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT5), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G176gat), .B(G204gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT68), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n540_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT69), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n550_), .A2(new_n560_), .A3(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT13), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n564_), .A3(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT70), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G29gat), .B(G36gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n571_), .A2(new_n573_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n568_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n569_), .B(new_n570_), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n572_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(KEYINPUT15), .A3(new_n574_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n577_), .A2(new_n546_), .A3(new_n580_), .A4(new_n547_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n574_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(new_n508_), .A3(new_n534_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT34), .Z(new_n585_));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n588_), .A2(KEYINPUT74), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(KEYINPUT74), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n585_), .A2(new_n586_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n581_), .A2(new_n583_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n581_), .A2(new_n583_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n587_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n581_), .A2(KEYINPUT75), .A3(new_n583_), .A4(new_n592_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G190gat), .B(G218gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT73), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT76), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n604_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n599_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n605_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n599_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n612_), .B(new_n613_), .C1(new_n608_), .C2(new_n599_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n614_), .A3(KEYINPUT77), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT77), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n616_), .B(KEYINPUT37), .C1(new_n607_), .C2(new_n609_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G15gat), .B(G22gat), .ZN(new_n619_));
  INV_X1    g418(.A(G1gat), .ZN(new_n620_));
  INV_X1    g419(.A(G8gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT14), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G1gat), .B(G8gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT78), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT79), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n526_), .B(new_n628_), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n626_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT16), .ZN(new_n633_));
  XOR2_X1   g432(.A(G183gat), .B(G211gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n630_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(KEYINPUT17), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n630_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n618_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n625_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n577_), .A2(new_n640_), .A3(new_n580_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n582_), .B2(new_n625_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n582_), .A2(new_n625_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n579_), .A3(new_n574_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n641_), .A2(new_n644_), .B1(new_n647_), .B2(new_n643_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G113gat), .B(G141gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G169gat), .B(G197gat), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n649_), .B(new_n650_), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n648_), .B(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR4_X1   g452(.A1(new_n490_), .A2(new_n567_), .A3(new_n639_), .A4(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT105), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(KEYINPUT105), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n657_), .A2(G1gat), .A3(new_n458_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT38), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(KEYINPUT38), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n609_), .B1(new_n599_), .B2(new_n611_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n490_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n566_), .B2(new_n653_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n566_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(KEYINPUT106), .A3(new_n652_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n662_), .A2(new_n638_), .A3(new_n664_), .A4(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G1gat), .B1(new_n667_), .B2(new_n458_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n659_), .A2(new_n660_), .A3(new_n668_), .ZN(G1324gat));
  OAI21_X1  g468(.A(G8gat), .B1(new_n667_), .B2(new_n332_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(KEYINPUT39), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(KEYINPUT39), .ZN(new_n672_));
  INV_X1    g471(.A(new_n332_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n621_), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n671_), .A2(new_n672_), .B1(new_n657_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  OAI221_X1 g477(.A(new_n676_), .B1(new_n657_), .B2(new_n674_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  INV_X1    g479(.A(new_n358_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G15gat), .B1(new_n667_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n683_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n681_), .A2(G15gat), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n684_), .A2(new_n685_), .B1(new_n657_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI221_X1 g488(.A(KEYINPUT108), .B1(new_n657_), .B2(new_n686_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1326gat));
  OAI21_X1  g490(.A(G22gat), .B1(new_n667_), .B2(new_n419_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n419_), .A2(G22gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n657_), .B2(new_n695_), .ZN(G1327gat));
  NOR2_X1   g495(.A1(new_n490_), .A2(new_n653_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n638_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n661_), .A2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n566_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n458_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G29gat), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n666_), .A2(new_n698_), .A3(new_n664_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n615_), .A2(new_n617_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n707_), .B(new_n708_), .C1(new_n483_), .C2(new_n489_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n488_), .B1(new_n487_), .B2(new_n358_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n464_), .A2(new_n481_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(KEYINPUT104), .A3(new_n681_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n713_), .A3(new_n459_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n707_), .B1(new_n714_), .B2(new_n708_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n706_), .B1(new_n710_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n706_), .C1(new_n710_), .C2(new_n715_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n703_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n704_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  NOR2_X1   g523(.A1(new_n332_), .A2(G36gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n702_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n726_), .B(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n719_), .A2(new_n673_), .A3(new_n720_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n719_), .A2(KEYINPUT111), .A3(new_n673_), .A4(new_n720_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G36gat), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n729_), .B(KEYINPUT46), .C1(new_n732_), .C2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n726_), .B(new_n727_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n733_), .A2(G36gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n730_), .A2(new_n731_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT113), .B(KEYINPUT46), .Z(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(G1329gat));
  NAND2_X1  g540(.A1(new_n358_), .A2(G43gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n701_), .A2(new_n681_), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n721_), .A2(new_n742_), .B1(G43gat), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g544(.A(G50gat), .B1(new_n702_), .B2(new_n462_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n462_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n722_), .B2(new_n747_), .ZN(G1331gat));
  NAND4_X1  g547(.A1(new_n662_), .A2(new_n653_), .A3(new_n567_), .A4(new_n638_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G57gat), .B1(new_n749_), .B2(new_n458_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n490_), .A2(new_n652_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n751_), .A2(new_n566_), .A3(new_n638_), .A4(new_n618_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n458_), .A2(G57gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1332gat));
  OAI21_X1  g553(.A(G64gat), .B1(new_n749_), .B2(new_n332_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT48), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n332_), .A2(G64gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n752_), .B2(new_n757_), .ZN(G1333gat));
  OAI21_X1  g557(.A(G71gat), .B1(new_n749_), .B2(new_n681_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT49), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n358_), .A2(new_n334_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n752_), .B2(new_n761_), .ZN(G1334gat));
  OAI21_X1  g561(.A(G78gat), .B1(new_n749_), .B2(new_n419_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT50), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n419_), .A2(G78gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n752_), .B2(new_n765_), .ZN(G1335gat));
  INV_X1    g565(.A(new_n567_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n699_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n751_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n492_), .A3(new_n703_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n665_), .A2(new_n652_), .A3(new_n638_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n490_), .B2(new_n618_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n709_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(new_n703_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n776_), .B2(new_n492_), .ZN(G1336gat));
  NAND3_X1  g576(.A1(new_n770_), .A2(new_n493_), .A3(new_n673_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n775_), .A2(new_n673_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n493_), .ZN(G1337gat));
  AOI21_X1  g579(.A(new_n511_), .B1(new_n775_), .B2(new_n358_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n358_), .A2(new_n503_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n769_), .A2(new_n782_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n781_), .A2(KEYINPUT114), .A3(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g584(.A1(new_n770_), .A2(new_n504_), .A3(new_n462_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n775_), .A2(new_n462_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(G106gat), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT52), .B(new_n504_), .C1(new_n775_), .C2(new_n462_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT53), .ZN(G1339gat));
  XOR2_X1   g591(.A(KEYINPUT118), .B(G113gat), .Z(new_n793_));
  NAND2_X1  g592(.A1(new_n652_), .A2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT119), .Z(new_n795_));
  NOR2_X1   g594(.A1(new_n673_), .A2(new_n462_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n358_), .A3(new_n703_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n651_), .B1(new_n647_), .B2(new_n642_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n641_), .A2(new_n645_), .A3(new_n643_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n648_), .A2(new_n651_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n558_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT116), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n558_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n544_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n549_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n543_), .A2(new_n548_), .A3(KEYINPUT55), .A4(new_n544_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n556_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n812_), .B(new_n555_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n805_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n805_), .B(KEYINPUT58), .C1(new_n811_), .C2(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n708_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n559_), .A2(new_n561_), .A3(new_n800_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n652_), .A2(new_n558_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n819_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n820_), .B(KEYINPUT115), .C1(new_n811_), .C2(new_n813_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n661_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n818_), .B1(new_n825_), .B2(KEYINPUT57), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n827_), .B(new_n661_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n698_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n638_), .A2(new_n653_), .ZN(new_n830_));
  OR4_X1    g629(.A1(KEYINPUT54), .A2(new_n708_), .A3(new_n566_), .A4(new_n830_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n566_), .A2(new_n830_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT54), .B1(new_n832_), .B2(new_n708_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n797_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n837_), .B(new_n797_), .C1(new_n829_), .C2(new_n834_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n795_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  AOI211_X1 g638(.A(KEYINPUT117), .B(G113gat), .C1(new_n835_), .C2(new_n652_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n829_), .A2(new_n834_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n797_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n652_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(G113gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n839_), .B1(new_n840_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n839_), .B(KEYINPUT120), .C1(new_n846_), .C2(new_n840_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1340gat));
  NOR2_X1   g650(.A1(new_n836_), .A2(new_n838_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852_), .B2(new_n767_), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n665_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n835_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n852_), .B2(new_n698_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n835_), .A2(new_n342_), .A3(new_n638_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1342gat));
  OAI21_X1  g659(.A(G134gat), .B1(new_n852_), .B2(new_n618_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n835_), .A2(new_n340_), .A3(new_n661_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n358_), .A2(new_n419_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(new_n673_), .A3(new_n458_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n842_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n653_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT121), .B(G141gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n867_), .A2(new_n767_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n369_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n867_), .A2(new_n698_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT122), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT123), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n873_), .B(new_n876_), .ZN(G1346gat));
  INV_X1    g676(.A(new_n867_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n878_), .A2(G162gat), .A3(new_n708_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G162gat), .B1(new_n878_), .B2(new_n661_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n881_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(G1347gat));
  AOI21_X1  g683(.A(new_n332_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n681_), .A2(new_n462_), .A3(new_n703_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n217_), .B1(new_n887_), .B2(new_n652_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n888_), .A2(KEYINPUT62), .ZN(new_n889_));
  INV_X1    g688(.A(new_n887_), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n890_), .A2(new_n300_), .A3(new_n653_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(KEYINPUT62), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n891_), .A3(new_n892_), .ZN(G1348gat));
  OAI21_X1  g692(.A(G176gat), .B1(new_n890_), .B2(new_n767_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n887_), .A2(new_n218_), .A3(new_n566_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1349gat));
  AOI21_X1  g695(.A(G183gat), .B1(new_n887_), .B2(new_n638_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n890_), .A2(new_n698_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n286_), .A2(new_n291_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n890_), .B2(new_n618_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n661_), .A2(new_n287_), .A3(new_n294_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n890_), .B2(new_n902_), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n865_), .A2(new_n703_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n332_), .B(new_n905_), .C1(new_n829_), .C2(new_n834_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n652_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g707(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT125), .B(G204gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n567_), .ZN(new_n911_));
  MUX2_X1   g710(.A(new_n909_), .B(new_n910_), .S(new_n911_), .Z(G1353gat));
  NAND2_X1  g711(.A1(new_n906_), .A2(new_n638_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT63), .B(G211gat), .Z(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n913_), .B2(new_n915_), .ZN(G1354gat));
  NAND3_X1  g715(.A1(new_n906_), .A2(G218gat), .A3(new_n708_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n885_), .A2(new_n918_), .A3(new_n661_), .A4(new_n904_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n254_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n906_), .B2(new_n661_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n917_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT127), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n924_), .B(new_n917_), .C1(new_n920_), .C2(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1355gat));
endmodule


