//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT10), .B(G99gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G92gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n208_), .A2(G85gat), .B1(KEYINPUT9), .B2(new_n209_), .ZN(new_n210_));
  AND3_X1   g009(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  OAI221_X1 g010(.A(new_n206_), .B1(G106gat), .B2(new_n207_), .C1(new_n210_), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n206_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT7), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n206_), .A2(new_n214_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G85gat), .B(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n213_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  AOI211_X1 g021(.A(KEYINPUT8), .B(new_n220_), .C1(new_n217_), .C2(new_n206_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n212_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G57gat), .B(G64gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n226_));
  XOR2_X1   g025(.A(G71gat), .B(G78gat), .Z(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n226_), .A2(new_n227_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n224_), .A2(new_n231_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT12), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT12), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n224_), .A2(new_n235_), .A3(new_n231_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n204_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n238_));
  INV_X1    g037(.A(new_n232_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n233_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n204_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G120gat), .B(G148gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT5), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G176gat), .B(G204gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n243_), .A2(new_n247_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n202_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(KEYINPUT13), .A3(new_n248_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT67), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT14), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT74), .B(G1gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(G8gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G15gat), .B(G22gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G1gat), .B(G8gat), .Z(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G231gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT76), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n266_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(new_n231_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G127gat), .B(G155gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT16), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G183gat), .B(G211gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n275_));
  OR3_X1    g074(.A1(new_n270_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n274_), .B(KEYINPUT17), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n270_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n270_), .B2(new_n278_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G43gat), .B(G50gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT68), .B(KEYINPUT15), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n224_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n283_), .B1(new_n224_), .B2(new_n288_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT71), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n286_), .B(new_n212_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G232gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT34), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT35), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT70), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n294_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT35), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n291_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G190gat), .B(G218gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G134gat), .B(G162gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT36), .ZN(new_n306_));
  INV_X1    g105(.A(new_n301_), .ZN(new_n307_));
  OAI221_X1 g106(.A(new_n297_), .B1(KEYINPUT71), .B2(new_n307_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n302_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT72), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n302_), .A2(new_n311_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n308_), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n305_), .B(KEYINPUT36), .Z(new_n314_));
  AOI22_X1  g113(.A1(new_n310_), .A2(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT37), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(KEYINPUT37), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n255_), .A2(new_n282_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT102), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT89), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT89), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(G155gat), .A3(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT1), .ZN(new_n329_));
  INV_X1    g128(.A(G155gat), .ZN(new_n330_));
  INV_X1    g129(.A(G162gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT88), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT88), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(G155gat), .B2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n325_), .A2(new_n327_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n329_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G141gat), .ZN(new_n340_));
  INV_X1    g139(.A(G148gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n335_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n339_), .A2(new_n344_), .B1(new_n345_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(G78gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G106gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n357_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G211gat), .B(G218gat), .Z(new_n364_));
  XOR2_X1   g163(.A(G197gat), .B(G204gat), .Z(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(KEYINPUT92), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G197gat), .B(G204gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT92), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT21), .B(new_n364_), .C1(new_n366_), .C2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT21), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n364_), .B1(new_n371_), .B2(new_n367_), .ZN(new_n372_));
  INV_X1    g171(.A(G197gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT21), .B(new_n374_), .C1(new_n365_), .C2(KEYINPUT91), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n370_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n363_), .A2(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n357_), .A2(new_n362_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n357_), .A2(new_n362_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(G71gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G99gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G43gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n391_), .B(new_n394_), .Z(new_n395_));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT23), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G183gat), .A3(G190gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n397_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT82), .B1(new_n398_), .B2(KEYINPUT23), .ZN(new_n403_));
  INV_X1    g202(.A(G183gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT80), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G183gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  OAI22_X1  g207(.A1(new_n402_), .A2(new_n403_), .B1(new_n408_), .B2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(G169gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT22), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT22), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(G176gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT81), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n409_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n422_));
  INV_X1    g221(.A(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT26), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT26), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G190gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT25), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n427_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n399_), .A2(new_n401_), .ZN(new_n432_));
  OR3_X1    g231(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n410_), .A2(new_n414_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT24), .A3(new_n416_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .A4(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n421_), .A2(new_n422_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n422_), .B1(new_n421_), .B2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n396_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n421_), .A2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT83), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n421_), .A2(new_n436_), .A3(new_n422_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(KEYINPUT30), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT86), .B1(new_n439_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n443_), .A3(KEYINPUT86), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n395_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n395_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G127gat), .B(G134gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G113gat), .B(G120gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n451_), .B(new_n452_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n450_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT31), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OR3_X1    g256(.A1(new_n447_), .A2(new_n449_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n457_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n386_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT19), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n424_), .B(new_n426_), .C1(new_n464_), .C2(new_n430_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n465_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n432_), .A2(KEYINPUT82), .ZN(new_n467_));
  INV_X1    g266(.A(new_n403_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n465_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n403_), .B1(new_n432_), .B2(KEYINPUT82), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT93), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n411_), .A2(new_n413_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n477_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n414_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n404_), .A2(new_n423_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n432_), .A2(new_n481_), .B1(G169gat), .B2(G176gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n475_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT20), .B(new_n463_), .C1(new_n484_), .C2(new_n377_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n370_), .A2(new_n376_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n484_), .B2(new_n377_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n441_), .A2(new_n442_), .A3(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n494_), .B2(new_n462_), .ZN(new_n495_));
  AOI211_X1 g294(.A(KEYINPUT95), .B(new_n463_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n489_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G8gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT18), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n437_), .A2(new_n438_), .A3(new_n377_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n471_), .A2(new_n474_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT20), .B1(new_n505_), .B2(new_n486_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n462_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT95), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n494_), .A2(new_n490_), .A3(new_n462_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(new_n489_), .A3(new_n501_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n503_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT27), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n466_), .A2(new_n469_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n486_), .A2(new_n483_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT20), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n462_), .B1(new_n517_), .B2(new_n487_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n462_), .B2(new_n494_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n513_), .B1(new_n519_), .B2(new_n502_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n511_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n460_), .A2(new_n514_), .A3(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G29gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G85gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT0), .B(G57gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n325_), .A2(new_n327_), .A3(new_n337_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n337_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n335_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n344_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n352_), .A2(new_n336_), .A3(new_n328_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n455_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n454_), .B(new_n533_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT4), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n455_), .B(new_n540_), .C1(new_n532_), .C2(new_n534_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n538_), .B(KEYINPUT97), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n451_), .A2(new_n452_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n451_), .A2(new_n452_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n450_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n453_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n536_), .B(KEYINPUT4), .C1(new_n549_), .C2(new_n353_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT96), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n535_), .A2(new_n552_), .A3(KEYINPUT4), .A4(new_n536_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n543_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n539_), .B1(new_n554_), .B2(KEYINPUT98), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n556_));
  AOI211_X1 g355(.A(new_n556_), .B(new_n543_), .C1(new_n551_), .C2(new_n553_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n527_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT100), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT100), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n560_), .B(new_n527_), .C1(new_n555_), .C2(new_n557_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n551_), .A2(new_n553_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n556_), .B1(new_n562_), .B2(new_n543_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n554_), .A2(KEYINPUT98), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n563_), .A2(new_n526_), .A3(new_n564_), .A4(new_n539_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n323_), .B1(new_n522_), .B2(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n512_), .A2(new_n513_), .B1(new_n511_), .B2(new_n520_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n566_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(KEYINPUT102), .A4(new_n460_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n526_), .B1(new_n537_), .B2(new_n542_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n541_), .A2(new_n538_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n572_), .B1(new_n562_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n503_), .A2(new_n511_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT33), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT99), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n565_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n565_), .A2(new_n577_), .A3(new_n576_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n519_), .A2(KEYINPUT32), .A3(new_n501_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n497_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n501_), .A2(KEYINPUT32), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n579_), .A2(new_n580_), .B1(new_n566_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT101), .B1(new_n585_), .B2(new_n386_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n501_), .B1(new_n510_), .B2(new_n489_), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n502_), .B(new_n488_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n555_), .A2(new_n557_), .A3(new_n527_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT33), .B1(new_n590_), .B2(KEYINPUT99), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n589_), .A2(new_n591_), .A3(new_n580_), .A4(new_n574_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n566_), .A2(new_n584_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n386_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n568_), .A2(new_n569_), .A3(new_n386_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n458_), .A2(new_n459_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n571_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n266_), .B(new_n286_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n264_), .A2(new_n265_), .A3(new_n288_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n266_), .B2(new_n286_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n602_), .A2(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT79), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G169gat), .B(G197gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n607_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n601_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n322_), .A2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT103), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT103), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n569_), .A2(new_n257_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n618_), .A2(KEYINPUT38), .A3(new_n619_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n601_), .A2(new_n315_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n254_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n612_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n281_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n569_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n623_), .A3(new_n629_), .ZN(G1324gat));
  NOR2_X1   g429(.A1(new_n568_), .A2(G8gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n616_), .A2(new_n617_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G8gat), .B1(new_n628_), .B2(new_n568_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n636_), .B(G8gat), .C1(new_n628_), .C2(new_n568_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n634_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n635_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n632_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n632_), .B(new_n641_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  OAI21_X1  g444(.A(G15gat), .B1(new_n628_), .B2(new_n600_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT41), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n615_), .A2(G15gat), .A3(new_n600_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1326gat));
  XNOR2_X1  g448(.A(new_n386_), .B(KEYINPUT106), .ZN(new_n650_));
  OAI21_X1  g449(.A(G22gat), .B1(new_n628_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n650_), .A2(G22gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n615_), .B2(new_n653_), .ZN(G1327gat));
  NAND2_X1  g453(.A1(new_n281_), .A2(new_n315_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n254_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n614_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT109), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n614_), .A2(new_n659_), .A3(new_n656_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(G29gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n566_), .A2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT110), .Z(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n597_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT101), .B(new_n386_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n600_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n567_), .A2(new_n570_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n321_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT107), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(KEYINPUT43), .C1(new_n601_), .C2(new_n321_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n671_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n626_), .A2(new_n282_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n678_), .A2(new_n680_), .A3(new_n569_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n665_), .B1(new_n681_), .B2(new_n662_), .ZN(G1328gat));
  OR2_X1    g481(.A1(new_n568_), .A2(KEYINPUT111), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n568_), .A2(KEYINPUT111), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(G36gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n658_), .A2(new_n660_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT45), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n658_), .A2(new_n690_), .A3(new_n660_), .A4(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n678_), .A2(new_n680_), .A3(new_n568_), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT46), .B(new_n692_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1329gat));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n677_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n677_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT43), .B(new_n321_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n601_), .B2(new_n321_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(KEYINPUT107), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n705_), .B2(new_n674_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n599_), .B(new_n701_), .C1(new_n706_), .C2(new_n679_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G43gat), .ZN(new_n708_));
  INV_X1    g507(.A(G43gat), .ZN(new_n709_));
  AND4_X1   g508(.A1(new_n709_), .A2(new_n658_), .A3(new_n599_), .A4(new_n660_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n700_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT47), .B(new_n710_), .C1(new_n707_), .C2(G43gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1330gat));
  INV_X1    g513(.A(G50gat), .ZN(new_n715_));
  INV_X1    g514(.A(new_n650_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n661_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n386_), .B(new_n701_), .C1(new_n706_), .C2(new_n679_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT112), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G50gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(KEYINPUT112), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1331gat));
  NOR2_X1   g521(.A1(new_n601_), .A2(new_n612_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(new_n254_), .A3(new_n282_), .A4(new_n321_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT113), .ZN(new_n725_));
  INV_X1    g524(.A(G57gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n566_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n255_), .A2(new_n612_), .A3(new_n281_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n624_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n569_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n725_), .A2(new_n733_), .A3(new_n685_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n729_), .B2(new_n685_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n735_), .A2(new_n736_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n725_), .A2(new_n388_), .A3(new_n599_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G71gat), .B1(new_n730_), .B2(new_n600_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT49), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT49), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(G1334gat));
  NAND3_X1  g543(.A1(new_n725_), .A2(new_n359_), .A3(new_n716_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G78gat), .B1(new_n730_), .B2(new_n650_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT50), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT50), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1335gat));
  NOR4_X1   g548(.A1(new_n255_), .A2(new_n601_), .A3(new_n612_), .A4(new_n655_), .ZN(new_n750_));
  INV_X1    g549(.A(G85gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n566_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n254_), .A2(new_n613_), .A3(new_n281_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n676_), .A2(KEYINPUT115), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n672_), .A2(new_n674_), .A3(new_n755_), .A4(new_n675_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n566_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n752_), .B1(new_n758_), .B2(new_n751_), .ZN(G1336gat));
  INV_X1    g558(.A(new_n568_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G92gat), .B1(new_n750_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n685_), .A2(new_n208_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT116), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n757_), .B2(new_n763_), .ZN(G1337gat));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  INV_X1    g564(.A(new_n207_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n750_), .A2(new_n599_), .A3(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n757_), .A2(new_n599_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n765_), .B(new_n767_), .C1(new_n768_), .C2(new_n390_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n390_), .B1(new_n757_), .B2(new_n599_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n767_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT51), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n750_), .A2(new_n361_), .A3(new_n386_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  INV_X1    g574(.A(new_n386_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n753_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n676_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n775_), .B1(new_n778_), .B2(G106gat), .ZN(new_n779_));
  AOI211_X1 g578(.A(KEYINPUT52), .B(new_n361_), .C1(new_n676_), .C2(new_n777_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n774_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g581(.A(G113gat), .ZN(new_n783_));
  INV_X1    g582(.A(new_n522_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n247_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n238_), .A2(new_n786_), .A3(new_n242_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n234_), .A2(new_n204_), .A3(new_n236_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(KEYINPUT55), .B2(new_n237_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n785_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  OR3_X1    g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n250_), .A2(new_n613_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n611_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n266_), .A2(new_n286_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n607_), .A2(new_n611_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n796_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n315_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT57), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n805_), .B(new_n315_), .C1(new_n796_), .C2(new_n801_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n790_), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n790_), .A2(KEYINPUT56), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n790_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT120), .B1(new_n790_), .B2(KEYINPUT56), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n808_), .A2(new_n811_), .A3(new_n812_), .A4(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n252_), .A2(new_n800_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n321_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n815_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n282_), .B1(new_n807_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n281_), .A2(new_n612_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n251_), .A2(new_n824_), .A3(new_n253_), .A4(KEYINPUT117), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n823_), .B1(new_n829_), .B2(new_n321_), .ZN(new_n830_));
  AOI211_X1 g629(.A(KEYINPUT54), .B(new_n819_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n566_), .B(new_n784_), .C1(new_n822_), .C2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n783_), .B1(new_n833_), .B2(new_n613_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT121), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n783_), .C1(new_n833_), .C2(new_n613_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n822_), .A2(new_n832_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(KEYINPUT59), .A3(new_n566_), .A4(new_n784_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n833_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n613_), .A2(new_n783_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n835_), .A2(new_n837_), .B1(new_n842_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g643(.A(new_n833_), .ZN(new_n845_));
  INV_X1    g644(.A(G120gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(KEYINPUT60), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n625_), .B2(KEYINPUT60), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(KEYINPUT122), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n845_), .B(new_n849_), .C1(KEYINPUT122), .C2(new_n848_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n255_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n846_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n845_), .B2(new_n282_), .ZN(new_n853_));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n282_), .B2(KEYINPUT123), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(KEYINPUT123), .B2(new_n854_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n842_), .B2(new_n856_), .ZN(G1342gat));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n845_), .A2(new_n858_), .A3(new_n315_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n321_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n858_), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n599_), .A2(new_n776_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n685_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n838_), .A2(new_n566_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n340_), .A3(new_n612_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G141gat), .B1(new_n865_), .B2(new_n613_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1344gat));
  INV_X1    g668(.A(new_n255_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n866_), .A2(new_n341_), .A3(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G148gat), .B1(new_n865_), .B2(new_n255_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1345gat));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  OR3_X1    g673(.A1(new_n865_), .A2(new_n281_), .A3(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n865_), .B2(new_n281_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1346gat));
  NOR2_X1   g676(.A1(new_n321_), .A2(new_n331_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT124), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n838_), .A2(new_n566_), .A3(new_n315_), .A4(new_n864_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n866_), .A2(new_n879_), .B1(new_n880_), .B2(new_n331_), .ZN(G1347gat));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n686_), .A2(new_n566_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n599_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n716_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n612_), .B(new_n885_), .C1(new_n822_), .C2(new_n832_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n886_), .B2(G169gat), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(new_n882_), .A3(G169gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(KEYINPUT62), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n478_), .A2(new_n479_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n886_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n887_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n890_), .A2(new_n894_), .ZN(G1348gat));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n254_), .B(new_n885_), .C1(new_n822_), .C2(new_n832_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(G176gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n897_), .A2(KEYINPUT126), .A3(new_n414_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n822_), .A2(new_n832_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n386_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n255_), .A2(new_n414_), .A3(new_n884_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n899_), .A2(new_n900_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NAND4_X1  g703(.A1(new_n902_), .A2(new_n599_), .A3(new_n282_), .A4(new_n883_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n408_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n901_), .A2(new_n716_), .A3(new_n884_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n281_), .A2(new_n430_), .A3(new_n464_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n905_), .A2(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n427_), .A3(new_n315_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n819_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(new_n423_), .ZN(G1351gat));
  NOR3_X1   g712(.A1(new_n686_), .A2(new_n566_), .A3(new_n863_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n901_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n612_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n870_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g719(.A(KEYINPUT63), .B(G211gat), .Z(new_n921_));
  AND3_X1   g720(.A1(new_n916_), .A2(new_n282_), .A3(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n282_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1354gat));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n916_), .A2(new_n926_), .A3(new_n315_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n916_), .A2(new_n819_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n929_), .B2(new_n926_), .ZN(G1355gat));
endmodule


