//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_;
  XNOR2_X1  g000(.A(KEYINPUT18), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT22), .B(G169gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT95), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n209_), .B2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT96), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(KEYINPUT96), .B(new_n207_), .C1(new_n209_), .C2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n217_), .B(new_n218_), .C1(G183gat), .C2(G190gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n213_), .A3(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n217_), .A2(new_n218_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT24), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n221_), .A2(new_n224_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n220_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G211gat), .B(G218gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G204gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n233_), .ZN(new_n238_));
  OAI211_X1 g037(.A(KEYINPUT21), .B(new_n237_), .C1(new_n238_), .C2(KEYINPUT88), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(KEYINPUT89), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n234_), .A2(KEYINPUT89), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n233_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n239_), .A2(new_n232_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT90), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n239_), .A2(KEYINPUT90), .A3(new_n232_), .A4(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n235_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n231_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT19), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT20), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT76), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT22), .B1(new_n254_), .B2(new_n225_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT22), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT76), .A3(G169gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n226_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT77), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n255_), .A2(KEYINPUT77), .A3(new_n226_), .A4(new_n257_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(new_n207_), .A3(new_n219_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n230_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n253_), .B1(new_n247_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n249_), .A2(new_n252_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT101), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n249_), .A2(KEYINPUT101), .A3(new_n252_), .A4(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n231_), .A2(KEYINPUT100), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT100), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n220_), .A2(new_n272_), .A3(new_n230_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n247_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n253_), .B1(new_n248_), .B2(new_n263_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n252_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n206_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n231_), .A2(new_n248_), .ZN(new_n278_));
  OAI211_X1 g077(.A(KEYINPUT20), .B(new_n252_), .C1(new_n247_), .C2(new_n264_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n249_), .A2(new_n265_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n251_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n283_), .A3(new_n205_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n277_), .A2(KEYINPUT27), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n252_), .B1(new_n249_), .B2(new_n265_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n206_), .B1(new_n286_), .B2(new_n280_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n287_), .A3(KEYINPUT97), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(new_n280_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT97), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n205_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n289_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n285_), .A2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT84), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT84), .ZN(new_n303_));
  OAI221_X1 g102(.A(new_n303_), .B1(new_n299_), .B2(new_n300_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n300_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT82), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT85), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n298_), .A2(new_n299_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322_));
  INV_X1    g121(.A(G113gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G120gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n322_), .B(G113gat), .ZN(new_n326_));
  INV_X1    g125(.A(G120gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n321_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n321_), .A2(new_n334_), .A3(new_n329_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n335_), .B(new_n336_), .C1(new_n330_), .C2(new_n334_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G85gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(G1gat), .B(G29gat), .Z(new_n341_));
  XOR2_X1   g140(.A(new_n340_), .B(new_n341_), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n333_), .A2(new_n337_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n294_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n321_), .A2(KEYINPUT29), .ZN(new_n348_));
  XOR2_X1   g147(.A(G22gat), .B(G50gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT28), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n348_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(KEYINPUT87), .Z(new_n353_));
  NOR2_X1   g152(.A1(new_n247_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n310_), .B2(new_n320_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(KEYINPUT86), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT86), .ZN(new_n358_));
  AOI211_X1 g157(.A(new_n358_), .B(new_n355_), .C1(new_n310_), .C2(new_n320_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n354_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT91), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n354_), .B(new_n362_), .C1(new_n357_), .C2(new_n359_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n352_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT92), .B(new_n364_), .C1(new_n356_), .C2(new_n247_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n356_), .B2(new_n247_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT92), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n361_), .A2(new_n363_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G78gat), .B(G106gat), .Z(new_n370_));
  AOI21_X1  g169(.A(new_n351_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT93), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n365_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n356_), .B(KEYINPUT86), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n362_), .B1(new_n375_), .B2(new_n354_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n363_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n374_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n370_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(KEYINPUT93), .A3(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n371_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n378_), .B1(KEYINPUT94), .B2(new_n370_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n369_), .A2(new_n383_), .A3(new_n379_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n351_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G71gat), .B(G99gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n262_), .A2(new_n387_), .A3(new_n230_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n262_), .B2(new_n230_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n263_), .A2(KEYINPUT30), .ZN(new_n391_));
  INV_X1    g190(.A(new_n386_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n262_), .A2(new_n387_), .A3(new_n230_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(G15gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G43gat), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n390_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT78), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n390_), .A2(new_n394_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n398_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n390_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT31), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n325_), .A2(new_n328_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n408_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n326_), .A2(new_n327_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n324_), .A2(G120gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT79), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n325_), .A2(new_n328_), .A3(new_n409_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT31), .A3(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n412_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n413_), .B1(new_n412_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n401_), .A2(new_n407_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n412_), .A2(new_n418_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n423_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n381_), .A2(new_n385_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n347_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n288_), .A2(new_n292_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT33), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n433_), .A2(KEYINPUT98), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n345_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n331_), .A2(new_n336_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n335_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n436_), .B(new_n342_), .C1(new_n437_), .C2(new_n336_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n345_), .A2(new_n434_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n432_), .A2(new_n435_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT32), .B(new_n205_), .C1(new_n270_), .C2(new_n276_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n290_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT99), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n290_), .A2(KEYINPUT99), .A3(new_n442_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n346_), .A2(new_n441_), .A3(new_n445_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n440_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n381_), .A2(new_n385_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n428_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n431_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G8gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G1gat), .A2(G8gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT14), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n452_), .B(KEYINPUT71), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n458_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G231gat), .A2(G233gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  XNOR2_X1  g264(.A(G71gat), .B(G78gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G57gat), .A2(G64gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G57gat), .A2(G64gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT11), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G57gat), .ZN(new_n472_));
  INV_X1    g271(.A(G64gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT11), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n468_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n467_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n466_), .B(KEYINPUT11), .C1(new_n470_), .C2(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n478_), .A3(KEYINPUT65), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT72), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n465_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT16), .B(G183gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G211gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(G127gat), .B(G155gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT17), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n479_), .B(KEYINPUT67), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n465_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT73), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n499_));
  INV_X1    g298(.A(G99gat), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n502_), .A2(new_n505_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT8), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n500_), .A2(KEYINPUT10), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n500_), .A2(KEYINPUT10), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n501_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n505_), .A2(new_n506_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n509_), .A2(KEYINPUT9), .A3(new_n510_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .A4(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n508_), .A2(KEYINPUT8), .A3(new_n511_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT64), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n514_), .A2(KEYINPUT64), .A3(new_n521_), .A4(new_n522_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G29gat), .B(G36gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G43gat), .ZN(new_n529_));
  INV_X1    g328(.A(G50gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G43gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n528_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(G50gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n527_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n534_), .A3(KEYINPUT15), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT15), .B1(new_n531_), .B2(new_n534_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n523_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n537_), .A2(new_n541_), .A3(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(G134gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G162gat), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(KEYINPUT36), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT69), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n555_), .B(KEYINPUT36), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n551_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n559_), .B(KEYINPUT70), .Z(new_n565_));
  OAI21_X1  g364(.A(new_n558_), .B1(new_n552_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT37), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n498_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n451_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n525_), .A2(new_n526_), .A3(new_n483_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n483_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n508_), .A2(KEYINPUT8), .A3(new_n511_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT8), .B1(new_n508_), .B2(new_n511_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT64), .B1(new_n577_), .B2(new_n521_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n526_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n574_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n571_), .B1(new_n577_), .B2(new_n521_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n492_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n572_), .A2(new_n573_), .A3(new_n580_), .A4(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT66), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n573_), .B1(new_n580_), .B2(new_n570_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n236_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(G176gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(KEYINPUT68), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT66), .ZN(new_n595_));
  AOI211_X1 g394(.A(new_n595_), .B(new_n573_), .C1(new_n580_), .C2(new_n570_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n587_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n585_), .B1(new_n583_), .B2(KEYINPUT66), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n593_), .B1(new_n599_), .B2(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n598_), .A2(KEYINPUT13), .A3(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G229gat), .A2(G233gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n463_), .A2(new_n534_), .A3(new_n531_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n529_), .A2(new_n530_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n533_), .A2(G50gat), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n460_), .B(new_n462_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n609_), .A2(new_n612_), .A3(KEYINPUT74), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT74), .B1(new_n609_), .B2(new_n612_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n608_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n463_), .ZN(new_n616_));
  OAI211_X1 g415(.A(KEYINPUT75), .B(new_n616_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT15), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n535_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n463_), .B1(new_n619_), .B2(new_n538_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT75), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n536_), .B2(new_n463_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n617_), .B(new_n607_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(new_n225_), .ZN(new_n626_));
  INV_X1    g425(.A(G197gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n628_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n615_), .A2(new_n623_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n606_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n569_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n346_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n635_), .A2(G1gat), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT102), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n638_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n633_), .B(KEYINPUT103), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n497_), .B1(new_n431_), .B2(new_n450_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n562_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n636_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n641_), .A3(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(new_n294_), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n635_), .A2(G8gat), .A3(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .A4(new_n294_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(G8gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G8gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT104), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n649_), .B(new_n656_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g458(.A(G15gat), .B1(new_n645_), .B2(new_n428_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT41), .Z(new_n661_));
  INV_X1    g460(.A(new_n428_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n396_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n635_), .B2(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n645_), .B2(new_n449_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT105), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n667_), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n635_), .A2(G22gat), .A3(new_n449_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(G1327gat));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n564_), .A2(new_n567_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n451_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n564_), .A2(new_n567_), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT43), .B(new_n675_), .C1(new_n431_), .C2(new_n450_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n498_), .B(new_n642_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n677_), .A2(new_n681_), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n674_), .A2(new_n676_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n498_), .A4(new_n642_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n346_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n683_), .A2(KEYINPUT108), .A3(new_n346_), .A4(new_n685_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(G29gat), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n644_), .B1(new_n431_), .B2(new_n450_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(new_n634_), .A3(new_n498_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n693_), .A2(G29gat), .A3(new_n636_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n648_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n685_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n697_), .A3(new_n294_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n696_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n682_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n681_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n294_), .B(new_n685_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1329gat));
  OAI21_X1  g508(.A(new_n532_), .B1(new_n693_), .B2(new_n428_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n683_), .A2(new_n662_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n685_), .A2(G43gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n710_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  OAI21_X1  g516(.A(new_n530_), .B1(new_n693_), .B2(new_n449_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n449_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n683_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n685_), .A2(G50gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT109), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n724_), .B(new_n718_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n606_), .A2(new_n632_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n569_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n472_), .B1(new_n728_), .B2(new_n636_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n498_), .ZN(new_n730_));
  AND4_X1   g529(.A1(new_n644_), .A2(new_n451_), .A3(new_n730_), .A4(new_n727_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(G57gat), .A3(new_n346_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n729_), .A2(new_n732_), .ZN(G1332gat));
  AOI21_X1  g532(.A(new_n473_), .B1(new_n731_), .B2(new_n294_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT48), .Z(new_n735_));
  INV_X1    g534(.A(new_n728_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n473_), .A3(new_n294_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n731_), .B2(new_n662_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT49), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n739_), .A3(new_n662_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n731_), .A2(new_n719_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G78gat), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT50), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n728_), .A2(G78gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n449_), .B2(new_n747_), .ZN(G1335gat));
  AND3_X1   g547(.A1(new_n691_), .A2(new_n498_), .A3(new_n727_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n346_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n684_), .A2(new_n498_), .A3(new_n727_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n636_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n752_), .B2(G85gat), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n751_), .B2(new_n648_), .ZN(new_n754_));
  INV_X1    g553(.A(G92gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n749_), .A2(new_n755_), .A3(new_n294_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT110), .ZN(G1337gat));
  OAI211_X1 g557(.A(new_n749_), .B(new_n662_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT111), .ZN(new_n760_));
  OAI21_X1  g559(.A(G99gat), .B1(new_n751_), .B2(new_n428_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n749_), .A2(new_n501_), .A3(new_n719_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n684_), .A2(new_n498_), .A3(new_n719_), .A4(new_n727_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g570(.A1(new_n294_), .A2(new_n636_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n430_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n497_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n617_), .B(new_n608_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n628_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n631_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n594_), .B1(new_n587_), .B2(new_n597_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n599_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT114), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n601_), .A2(new_n784_), .A3(new_n779_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n527_), .A2(new_n574_), .B1(new_n581_), .B2(new_n492_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n572_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n573_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n583_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n787_), .A2(KEYINPUT55), .A3(new_n573_), .A4(new_n572_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n788_), .A2(KEYINPUT112), .A3(new_n789_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n792_), .A2(new_n794_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n591_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n591_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(KEYINPUT113), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n797_), .A2(new_n803_), .A3(KEYINPUT56), .A4(new_n591_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n587_), .A2(new_n592_), .A3(new_n597_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(new_n632_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n786_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n807_), .B2(new_n562_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n784_), .B1(new_n601_), .B2(new_n779_), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT114), .B(new_n778_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n591_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n591_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n803_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n804_), .A2(new_n632_), .A3(new_n805_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n812_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n644_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n808_), .A2(new_n809_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(KEYINPUT57), .A3(new_n644_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n805_), .B(new_n779_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n800_), .A2(new_n801_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(KEYINPUT58), .A3(new_n805_), .A4(new_n779_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n673_), .A2(new_n824_), .A3(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n821_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n774_), .B1(new_n820_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n632_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n568_), .A2(new_n606_), .A3(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT54), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n773_), .B1(new_n829_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n632_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n821_), .A2(new_n827_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n806_), .A2(new_n802_), .ZN(new_n838_));
  AOI211_X1 g637(.A(KEYINPUT115), .B(new_n562_), .C1(new_n838_), .C2(new_n812_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n818_), .B1(new_n817_), .B2(new_n644_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n837_), .B1(new_n841_), .B2(new_n809_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT117), .B1(new_n842_), .B2(new_n730_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n820_), .A2(new_n828_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n498_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n832_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n773_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n834_), .A2(KEYINPUT59), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n851_), .A2(new_n632_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n836_), .B1(new_n853_), .B2(G113gat), .ZN(G1340gat));
  AOI21_X1  g653(.A(new_n845_), .B1(new_n844_), .B2(new_n498_), .ZN(new_n855_));
  AOI211_X1 g654(.A(KEYINPUT117), .B(new_n730_), .C1(new_n820_), .C2(new_n828_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n833_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n605_), .B(new_n852_), .C1(new_n857_), .C2(new_n849_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n851_), .A2(KEYINPUT118), .A3(new_n605_), .A4(new_n852_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(G120gat), .A3(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n327_), .B1(new_n606_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n835_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n327_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1341gat));
  AOI21_X1  g664(.A(G127gat), .B1(new_n835_), .B2(new_n730_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n851_), .A2(new_n852_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n774_), .A2(G127gat), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT119), .Z(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n867_), .B2(new_n869_), .ZN(G1342gat));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871_));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n675_), .A2(new_n872_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n851_), .A2(new_n852_), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n834_), .B2(new_n644_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT120), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n872_), .C1(new_n834_), .C2(new_n644_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n871_), .B1(new_n874_), .B2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n851_), .A2(new_n852_), .A3(new_n873_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n881_), .A2(KEYINPUT121), .A3(new_n878_), .A4(new_n876_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1343gat));
  NOR2_X1   g682(.A1(new_n829_), .A2(new_n833_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n429_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(KEYINPUT122), .A3(new_n772_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n832_), .B1(new_n842_), .B2(new_n774_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(new_n429_), .A3(new_n772_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n830_), .B1(new_n887_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(G141gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1344gat));
  AOI21_X1  g693(.A(new_n606_), .B1(new_n887_), .B2(new_n891_), .ZN(new_n895_));
  INV_X1    g694(.A(G148gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1345gat));
  AOI21_X1  g696(.A(new_n498_), .B1(new_n887_), .B2(new_n891_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n898_), .B(new_n900_), .ZN(G1346gat));
  NAND2_X1  g700(.A1(new_n887_), .A2(new_n891_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n562_), .ZN(new_n903_));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n887_), .B2(new_n891_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n903_), .A2(new_n904_), .B1(new_n905_), .B2(new_n673_), .ZN(G1347gat));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n346_), .B1(new_n285_), .B2(new_n293_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n662_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n910_), .A2(KEYINPUT123), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(KEYINPUT123), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n830_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n913_), .A2(KEYINPUT124), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(KEYINPUT124), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n719_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n847_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n908_), .B1(new_n917_), .B2(G169gat), .ZN(new_n918_));
  AOI211_X1 g717(.A(KEYINPUT125), .B(new_n225_), .C1(new_n847_), .C2(new_n916_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n907_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n914_), .A2(new_n915_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n449_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n855_), .A2(new_n856_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n832_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT125), .B1(new_n924_), .B2(new_n225_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n917_), .A2(new_n908_), .A3(G169gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n925_), .A2(KEYINPUT62), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n719_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n847_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT126), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n847_), .A2(new_n931_), .A3(new_n928_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n830_), .A2(new_n209_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT127), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(new_n932_), .A3(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n920_), .A2(new_n927_), .A3(new_n935_), .ZN(G1348gat));
  NAND3_X1  g735(.A1(new_n930_), .A2(new_n605_), .A3(new_n932_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n888_), .A2(new_n928_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n606_), .A2(new_n226_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n937_), .A2(new_n226_), .B1(new_n938_), .B2(new_n939_), .ZN(G1349gat));
  AOI21_X1  g739(.A(G183gat), .B1(new_n938_), .B2(new_n730_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n930_), .A2(new_n932_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n497_), .A2(new_n222_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n941_), .B1(new_n942_), .B2(new_n943_), .ZN(G1350gat));
  NAND4_X1  g743(.A1(new_n930_), .A2(new_n562_), .A3(new_n223_), .A4(new_n932_), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n930_), .A2(new_n673_), .A3(new_n932_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n216_), .ZN(G1351gat));
  NAND2_X1  g746(.A1(new_n886_), .A2(new_n909_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n830_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(new_n627_), .ZN(G1352gat));
  NOR2_X1   g749(.A1(new_n948_), .A2(new_n606_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(new_n236_), .ZN(G1353gat));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  AND2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  NOR4_X1   g753(.A1(new_n948_), .A2(new_n497_), .A3(new_n953_), .A4(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n948_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n774_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n957_), .B2(new_n953_), .ZN(G1354gat));
  INV_X1    g757(.A(G218gat), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n948_), .A2(new_n959_), .A3(new_n675_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n956_), .A2(new_n562_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n959_), .B2(new_n961_), .ZN(G1355gat));
endmodule


