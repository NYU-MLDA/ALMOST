//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT86), .A3(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n206_));
  OAI21_X1  g005(.A(G169gat), .B1(new_n206_), .B2(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n205_), .A2(KEYINPUT87), .A3(new_n207_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n204_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n223_));
  OR3_X1    g022(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n215_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT25), .B(G183gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  OAI211_X1 g027(.A(KEYINPUT85), .B(G190gat), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT85), .A2(G190gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT84), .A3(KEYINPUT26), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n227_), .B1(new_n228_), .B2(G190gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n219_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G71gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G15gat), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT88), .B(G113gat), .ZN(new_n247_));
  INV_X1    g046(.A(G120gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT31), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n245_), .B1(new_n246_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n246_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n243_), .A2(new_n257_), .A3(new_n244_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  AND2_X1   g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n260_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(KEYINPUT1), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n260_), .B(KEYINPUT3), .Z(new_n269_));
  XOR2_X1   g068(.A(new_n267_), .B(KEYINPUT2), .Z(new_n270_));
  OAI21_X1  g069(.A(new_n263_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n254_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n268_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(KEYINPUT4), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT101), .B1(new_n274_), .B2(KEYINPUT4), .ZN(new_n276_));
  INV_X1    g075(.A(new_n254_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT101), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .A4(new_n273_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n272_), .A2(new_n274_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT0), .B(G57gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G85gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(G1gat), .B(G29gat), .Z(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n284_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n259_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT91), .ZN(new_n298_));
  INV_X1    g097(.A(G197gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(G204gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT92), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(G197gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n300_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT93), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT21), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n306_), .B2(KEYINPUT21), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G211gat), .A2(G218gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G211gat), .A2(G218gat), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT94), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT94), .ZN(new_n314_));
  OR2_X1    g113(.A1(G211gat), .A2(G218gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n299_), .A2(G204gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n302_), .A2(G197gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n313_), .A2(new_n316_), .B1(KEYINPUT21), .B2(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n308_), .A2(new_n309_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT94), .B1(new_n311_), .B2(new_n312_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n314_), .A3(new_n310_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT21), .A4(new_n319_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n226_), .A2(new_n327_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n215_), .A2(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n203_), .A2(new_n204_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n225_), .A2(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT95), .B1(new_n321_), .B2(new_n325_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n306_), .A2(KEYINPUT21), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n334_));
  INV_X1    g133(.A(new_n319_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n335_), .A2(new_n336_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT21), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n324_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n332_), .A2(new_n341_), .ZN(new_n342_));
  OAI221_X1 g141(.A(KEYINPUT20), .B1(new_n326_), .B2(new_n331_), .C1(new_n342_), .C2(new_n235_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT98), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n339_), .A2(new_n324_), .A3(new_n331_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT97), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT97), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n339_), .A2(new_n351_), .A3(new_n324_), .A4(new_n331_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n345_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n341_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n340_), .B1(new_n339_), .B2(new_n324_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n235_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AND4_X1   g156(.A1(new_n347_), .A2(new_n353_), .A3(new_n354_), .A4(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n345_), .B1(new_n342_), .B2(new_n235_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n347_), .B1(new_n359_), .B2(new_n353_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n346_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G8gat), .B(G36gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n346_), .B(new_n368_), .C1(new_n358_), .C2(new_n360_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(KEYINPUT100), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT100), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(new_n372_), .A3(new_n366_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n343_), .A2(new_n354_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n357_), .A2(KEYINPUT20), .A3(new_n345_), .A4(new_n349_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n366_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n369_), .A2(KEYINPUT27), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT96), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n355_), .A2(new_n356_), .ZN(new_n387_));
  AND2_X1   g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n326_), .B2(new_n389_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n390_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n395_));
  OR3_X1    g194(.A1(new_n386_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n384_), .A2(new_n385_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n397_), .B(new_n386_), .C1(new_n395_), .C2(new_n394_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n297_), .A2(new_n379_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n353_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT98), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n359_), .A2(new_n347_), .A3(new_n353_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n346_), .A3(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n375_), .A2(KEYINPUT32), .A3(new_n368_), .A4(new_n376_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n295_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n370_), .A2(new_n373_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n285_), .A2(new_n283_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n291_), .B(new_n413_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n291_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(KEYINPUT33), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT102), .B1(new_n293_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n419_), .A3(KEYINPUT33), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n416_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n411_), .B1(new_n412_), .B2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n259_), .B1(new_n422_), .B2(new_n399_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT103), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n400_), .B1(new_n379_), .B2(new_n295_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n402_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT67), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT66), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT7), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n432_), .A2(new_n433_), .B1(new_n237_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n237_), .A3(new_n434_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n429_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G99gat), .A2(G106gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT6), .ZN(new_n440_));
  INV_X1    g239(.A(new_n433_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n442_));
  OAI22_X1  g241(.A1(new_n441_), .A2(new_n442_), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT67), .A3(new_n436_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G85gat), .B(G92gat), .Z(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(KEYINPUT8), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n443_), .A3(new_n436_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n446_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G85gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n452_), .A2(G85gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(G92gat), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(KEYINPUT10), .B(G99gat), .Z(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT64), .B(G106gat), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n446_), .A2(KEYINPUT9), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n456_), .A2(new_n459_), .A3(new_n460_), .A4(new_n440_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G57gat), .B(G64gat), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n464_));
  XOR2_X1   g263(.A(G71gat), .B(G78gat), .Z(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n464_), .A2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n447_), .A2(new_n451_), .A3(new_n461_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G230gat), .A2(G233gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT68), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n447_), .A2(new_n451_), .A3(new_n461_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n468_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(KEYINPUT12), .A3(new_n474_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT68), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n469_), .A2(new_n479_), .A3(new_n470_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n472_), .A2(new_n477_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n469_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(G230gat), .A3(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT69), .B(G204gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G120gat), .B(G148gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT5), .B(G176gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n481_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n488_), .B(KEYINPUT70), .Z(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n492_));
  OR3_X1    g291(.A1(new_n490_), .A2(new_n492_), .A3(KEYINPUT13), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT13), .B1(new_n490_), .B2(new_n492_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498_));
  INV_X1    g297(.A(G29gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT71), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT71), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G29gat), .ZN(new_n502_));
  INV_X1    g301(.A(G36gat), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n500_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n501_), .A2(G29gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n499_), .A2(KEYINPUT71), .ZN(new_n508_));
  OAI21_X1  g307(.A(G36gat), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G43gat), .B(G50gat), .Z(new_n510_));
  NAND3_X1  g309(.A1(new_n500_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n506_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G1gat), .A2(G8gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT14), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT78), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT78), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n518_), .A3(KEYINPUT14), .ZN(new_n519_));
  INV_X1    g318(.A(G15gat), .ZN(new_n520_));
  INV_X1    g319(.A(G22gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G15gat), .A2(G22gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n517_), .A2(new_n519_), .A3(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G1gat), .B(G8gat), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(KEYINPUT78), .A2(new_n516_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n526_), .A3(new_n519_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n514_), .A2(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n504_), .A2(new_n505_), .A3(new_n498_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n510_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n528_), .B(new_n530_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT82), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n526_), .B1(new_n529_), .B2(new_n519_), .ZN(new_n539_));
  AND4_X1   g338(.A1(new_n526_), .A2(new_n517_), .A3(new_n519_), .A4(new_n524_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n512_), .B(new_n506_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n535_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT81), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n535_), .A3(KEYINPUT81), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(G229gat), .A3(G233gat), .A4(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(new_n220_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n299_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n538_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n538_), .B2(new_n546_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n497_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(KEYINPUT83), .A3(new_n551_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n496_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n447_), .A2(new_n513_), .A3(new_n451_), .A4(new_n461_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT72), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n473_), .A2(new_n514_), .B1(new_n562_), .B2(new_n561_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n569_), .ZN(new_n571_));
  AND4_X1   g370(.A1(new_n564_), .A2(new_n570_), .A3(new_n567_), .A4(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT76), .B1(new_n568_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(G134gat), .ZN(new_n575_));
  INV_X1    g374(.A(G162gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT36), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT73), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n570_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n563_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n566_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n573_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n581_), .A2(new_n582_), .A3(new_n588_), .A4(new_n577_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n573_), .A2(KEYINPUT77), .A3(new_n579_), .A4(new_n584_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT37), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT74), .B(new_n579_), .C1(new_n568_), .C2(new_n572_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n581_), .A2(new_n582_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT74), .B1(new_n595_), .B2(new_n579_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT37), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT75), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT75), .B(KEYINPUT37), .C1(new_n594_), .C2(new_n596_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n591_), .A2(new_n592_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n531_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n468_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n604_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT80), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n610_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n604_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n601_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n428_), .A2(new_n558_), .A3(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(KEYINPUT104), .ZN(new_n620_));
  INV_X1    g419(.A(G1gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(KEYINPUT104), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n295_), .A4(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(KEYINPUT105), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(KEYINPUT105), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n202_), .B1(new_n626_), .B2(KEYINPUT38), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n379_), .A2(new_n400_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n369_), .A2(KEYINPUT100), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n368_), .B1(new_n406_), .B2(new_n346_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n373_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n421_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n399_), .A3(new_n410_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n259_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n400_), .A2(new_n295_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .A4(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT103), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n401_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(new_n591_), .A3(new_n617_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n558_), .B(KEYINPUT106), .Z(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n621_), .B1(new_n643_), .B2(new_n295_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n626_), .B2(KEYINPUT38), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT107), .B(new_n646_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n627_), .A2(new_n645_), .A3(new_n647_), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n620_), .A2(new_n622_), .ZN(new_n649_));
  INV_X1    g448(.A(G8gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n379_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n379_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(G8gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n652_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  AOI21_X1  g458(.A(new_n520_), .B1(new_n643_), .B2(new_n259_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT41), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n649_), .A2(new_n520_), .A3(new_n259_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  AOI21_X1  g462(.A(new_n521_), .B1(new_n643_), .B2(new_n400_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT42), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n649_), .A2(new_n521_), .A3(new_n400_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1327gat));
  NAND2_X1  g466(.A1(new_n642_), .A2(new_n617_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n599_), .A2(new_n600_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(KEYINPUT37), .B2(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n640_), .A2(KEYINPUT43), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n428_), .B2(new_n601_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n669_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT44), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n640_), .B2(new_n672_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n428_), .A2(new_n674_), .A3(new_n601_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n668_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n681_), .A2(KEYINPUT108), .A3(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n296_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n640_), .A2(new_n671_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n617_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n496_), .A2(new_n557_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n499_), .A3(new_n295_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n691_), .ZN(G1328gat));
  OAI21_X1  g491(.A(new_n379_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G36gat), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(new_n379_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n428_), .A2(new_n591_), .A3(new_n688_), .A4(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT109), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .A4(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n695_), .A2(new_n696_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n676_), .A2(new_n677_), .A3(KEYINPUT44), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n682_), .B1(new_n681_), .B2(KEYINPUT108), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n503_), .B1(new_n707_), .B2(new_n379_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n700_), .B(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n703_), .B(new_n704_), .C1(new_n708_), .C2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n702_), .A2(new_n711_), .ZN(G1329gat));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713_));
  OAI21_X1  g512(.A(G43gat), .B1(new_n684_), .B2(new_n635_), .ZN(new_n714_));
  INV_X1    g513(.A(G43gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n690_), .A2(new_n715_), .A3(new_n259_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n635_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n713_), .B(new_n716_), .C1(new_n718_), .C2(new_n715_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n684_), .B2(new_n399_), .ZN(new_n722_));
  OR3_X1    g521(.A1(new_n689_), .A2(G50gat), .A3(new_n399_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1331gat));
  INV_X1    g523(.A(new_n557_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n495_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n428_), .A2(new_n618_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n295_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n641_), .A2(new_n726_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n296_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n731_), .B2(G57gat), .ZN(G1332gat));
  OAI21_X1  g531(.A(G64gat), .B1(new_n730_), .B2(new_n697_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT48), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n697_), .A2(G64gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n727_), .B2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n730_), .B2(new_n635_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n635_), .A2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n727_), .B2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n730_), .B2(new_n399_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n399_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n727_), .B2(new_n743_), .ZN(G1335gat));
  NOR3_X1   g543(.A1(new_n495_), .A2(new_n687_), .A3(new_n725_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n686_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n295_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n745_), .B(KEYINPUT111), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT112), .Z(new_n751_));
  INV_X1    g550(.A(new_n455_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n296_), .B2(new_n453_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n747_), .B1(new_n751_), .B2(new_n753_), .ZN(G1336gat));
  INV_X1    g553(.A(G92gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n746_), .A2(new_n755_), .A3(new_n379_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n751_), .A2(new_n379_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n755_), .ZN(G1337gat));
  AND3_X1   g557(.A1(new_n746_), .A2(new_n457_), .A3(new_n259_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n237_), .B1(new_n750_), .B2(new_n259_), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n759_), .A2(new_n760_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n761_));
  NAND2_X1  g560(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n746_), .A2(new_n458_), .A3(new_n400_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n750_), .A2(new_n400_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G106gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT52), .B(new_n434_), .C1(new_n750_), .C2(new_n400_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n481_), .A2(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n473_), .A2(KEYINPUT12), .A3(new_n474_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT12), .B1(new_n473_), .B2(new_n474_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(KEYINPUT55), .A3(new_n472_), .A4(new_n480_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n477_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(G230gat), .A3(G233gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n491_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(KEYINPUT56), .A3(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n544_), .A2(new_n545_), .A3(new_n537_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n549_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n788_), .B2(new_n549_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n537_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n532_), .A2(new_n535_), .A3(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n787_), .B1(new_n794_), .B2(new_n552_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n549_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT115), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(new_n789_), .A3(new_n549_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT116), .B(new_n551_), .C1(new_n799_), .C2(new_n793_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT117), .B1(new_n801_), .B2(new_n489_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n490_), .C1(new_n795_), .C2(new_n800_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n786_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n786_), .B(KEYINPUT58), .C1(new_n802_), .C2(new_n804_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n601_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n554_), .A2(new_n556_), .A3(new_n489_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n490_), .A2(new_n492_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n800_), .B2(new_n795_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n671_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n671_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT118), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n809_), .A2(new_n821_), .A3(new_n818_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n617_), .A3(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n496_), .A2(new_n725_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n618_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT54), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n672_), .A2(new_n827_), .A3(new_n687_), .A4(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT114), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n618_), .A2(new_n830_), .A3(new_n827_), .A4(new_n824_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n823_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n379_), .A2(new_n400_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n295_), .A3(new_n259_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n771_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT119), .B(new_n835_), .C1(new_n823_), .C2(new_n832_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n725_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n835_), .B1(new_n823_), .B2(new_n832_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n819_), .A2(new_n617_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n832_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n842_), .A3(new_n836_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n725_), .A2(G113gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT120), .Z(new_n849_));
  AOI21_X1  g648(.A(new_n840_), .B1(new_n847_), .B2(new_n849_), .ZN(G1340gat));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n496_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(KEYINPUT121), .A3(new_n496_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(G120gat), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n248_), .B1(new_n495_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n839_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n248_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n847_), .A2(G127gat), .A3(new_n687_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n687_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n860_));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n860_), .A2(KEYINPUT122), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT122), .B1(new_n860_), .B2(new_n861_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n859_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT123), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n859_), .B(new_n866_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1342gat));
  AOI21_X1  g667(.A(G134gat), .B1(new_n839_), .B2(new_n591_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n847_), .A2(G134gat), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n871_), .B2(new_n601_), .ZN(G1343gat));
  AOI21_X1  g671(.A(new_n636_), .B1(new_n823_), .B2(new_n832_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n379_), .A2(new_n259_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n725_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n875_), .A2(new_n495_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT124), .B(G148gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1345gat));
  NOR2_X1   g680(.A1(new_n875_), .A2(new_n617_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT61), .B(G155gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  NOR3_X1   g683(.A1(new_n875_), .A2(new_n576_), .A3(new_n672_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n876_), .A2(new_n591_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n576_), .B2(new_n886_), .ZN(G1347gat));
  NOR3_X1   g686(.A1(new_n697_), .A2(new_n297_), .A3(new_n400_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n845_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n557_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G169gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT62), .ZN(new_n893_));
  INV_X1    g692(.A(new_n203_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n891_), .ZN(G1348gat));
  INV_X1    g694(.A(new_n889_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G176gat), .B1(new_n896_), .B2(new_n496_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n204_), .B(new_n495_), .C1(new_n823_), .C2(new_n832_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n888_), .B2(new_n898_), .ZN(G1349gat));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n687_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n226_), .ZN(new_n901_));
  INV_X1    g700(.A(G183gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(KEYINPUT125), .B2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(KEYINPUT125), .B2(new_n901_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n889_), .B2(new_n672_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n591_), .A2(new_n327_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT126), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n889_), .B2(new_n908_), .ZN(G1351gat));
  NOR3_X1   g708(.A1(new_n628_), .A2(new_n295_), .A3(new_n259_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n833_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n725_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n299_), .A2(KEYINPUT127), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n299_), .A2(KEYINPUT127), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n915_), .ZN(G1352gat));
  NOR2_X1   g716(.A1(new_n911_), .A2(new_n495_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n302_), .ZN(G1353gat));
  NAND2_X1  g718(.A1(new_n912_), .A2(new_n687_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n920_), .B2(new_n921_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n911_), .A2(new_n925_), .A3(new_n672_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n912_), .A2(new_n591_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(G1355gat));
endmodule


