//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_,
    new_n977_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  XOR2_X1   g001(.A(G120gat), .B(G148gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G204gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT5), .B(G176gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT68), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n212_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(G85gat), .A4(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT65), .B1(new_n219_), .B2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n220_), .A2(new_n221_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n231_), .A2(new_n215_), .A3(new_n216_), .A4(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n229_), .A2(new_n230_), .A3(new_n212_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n210_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n238_), .A2(new_n225_), .A3(new_n226_), .A4(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n217_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT8), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT8), .B1(new_n240_), .B2(new_n241_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n235_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G57gat), .B(G64gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT11), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n248_));
  INV_X1    g047(.A(G57gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(G64gat), .ZN(new_n250_));
  INV_X1    g049(.A(G64gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(G57gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n248_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G71gat), .B(G78gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n247_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n246_), .A2(new_n254_), .A3(KEYINPUT11), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n208_), .B1(new_n245_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT12), .ZN(new_n262_));
  AOI211_X1 g061(.A(new_n258_), .B(new_n262_), .C1(new_n235_), .C2(new_n244_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n235_), .A2(new_n244_), .A3(new_n258_), .ZN(new_n265_));
  INV_X1    g064(.A(G230gat), .ZN(new_n266_));
  INV_X1    g065(.A(G233gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n235_), .A2(new_n244_), .A3(KEYINPUT66), .A4(new_n258_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n258_), .B1(new_n235_), .B2(new_n244_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n268_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n207_), .B1(new_n271_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n271_), .A2(new_n277_), .A3(new_n207_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT13), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT13), .B1(new_n279_), .B2(new_n280_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n202_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n281_), .A3(KEYINPUT69), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G29gat), .B(G36gat), .Z(new_n289_));
  XOR2_X1   g088(.A(G43gat), .B(G50gat), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G29gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G43gat), .B(G50gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT75), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n291_), .A2(KEYINPUT75), .A3(new_n294_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G1gat), .A2(G8gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT14), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G15gat), .A2(G22gat), .ZN(new_n301_));
  AND2_X1   g100(.A1(G15gat), .A2(G22gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT73), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT73), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G1gat), .B(G8gat), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n307_), .A3(new_n305_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n298_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n310_), .B(new_n309_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n291_), .A2(new_n294_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT15), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n291_), .A2(KEYINPUT15), .A3(new_n294_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n311_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G113gat), .B(G141gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G169gat), .ZN(new_n326_));
  INV_X1    g125(.A(G197gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n317_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n317_), .A2(new_n324_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n328_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n288_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G211gat), .B(G218gat), .Z(new_n339_));
  INV_X1    g138(.A(KEYINPUT21), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G197gat), .B(G204gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT21), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n342_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(KEYINPUT21), .A3(new_n343_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349_));
  OR2_X1    g148(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(G183gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n349_), .B1(new_n353_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n360_), .A2(KEYINPUT79), .A3(new_n356_), .A4(new_n357_), .ZN(new_n361_));
  INV_X1    g160(.A(G169gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT22), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G169gat), .ZN(new_n365_));
  INV_X1    g164(.A(G176gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(KEYINPUT78), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n367_), .A2(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n359_), .A2(new_n361_), .A3(new_n368_), .A4(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n350_), .A2(KEYINPUT26), .A3(new_n352_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT25), .B(G183gat), .ZN(new_n372_));
  INV_X1    g171(.A(G190gat), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n371_), .B(new_n372_), .C1(KEYINPUT26), .C2(new_n373_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n358_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT24), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n374_), .B(new_n376_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n348_), .A2(new_n370_), .A3(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n356_), .B(new_n357_), .C1(G183gat), .C2(G190gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n377_), .A3(new_n367_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n372_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n376_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n378_), .A2(KEYINPUT91), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT91), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n377_), .B2(KEYINPUT24), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n388_), .A2(new_n379_), .A3(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT92), .B1(new_n387_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n390_), .A2(new_n379_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(KEYINPUT91), .B2(new_n378_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT92), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n376_), .A4(new_n386_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n384_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n381_), .B(KEYINPUT20), .C1(new_n397_), .C2(new_n348_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n399_), .B(KEYINPUT89), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT90), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n400_), .A2(KEYINPUT19), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(KEYINPUT19), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT20), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n392_), .A2(new_n396_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n345_), .A2(new_n383_), .A3(new_n347_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n370_), .A2(new_n380_), .B1(new_n347_), .B2(new_n345_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n398_), .A2(new_n402_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT32), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G64gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(new_n214_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n412_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT97), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(new_n413_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n387_), .A2(new_n391_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT20), .B1(new_n407_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n401_), .B1(new_n410_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n419_), .A2(new_n420_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G57gat), .B(G85gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n436_), .B2(KEYINPUT84), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n438_), .A2(G141gat), .A3(G148gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n434_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(KEYINPUT84), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n438_), .B1(G141gat), .B2(G148gat), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(KEYINPUT85), .A3(new_n442_), .A4(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n447_), .B(new_n448_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G141gat), .A2(G148gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT82), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(G141gat), .A3(G148gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT2), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n444_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n457_), .A2(KEYINPUT1), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n457_), .B1(new_n459_), .B2(KEYINPUT1), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n463_), .B1(new_n464_), .B2(KEYINPUT83), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n466_), .B(new_n457_), .C1(new_n459_), .C2(KEYINPUT1), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n451_), .A2(new_n453_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(new_n436_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G127gat), .B(G134gat), .Z(new_n472_));
  XOR2_X1   g271(.A(G113gat), .B(G120gat), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G127gat), .B(G134gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G113gat), .B(G120gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n462_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT80), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n480_), .A3(new_n477_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(new_n476_), .A3(KEYINPUT80), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n460_), .B1(new_n444_), .B2(new_n455_), .ZN(new_n484_));
  AOI211_X1 g283(.A(new_n436_), .B(new_n469_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n433_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n462_), .A2(new_n471_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT4), .B1(new_n488_), .B2(new_n483_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n487_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n479_), .A2(new_n486_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n490_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n432_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(KEYINPUT4), .ZN(new_n496_));
  INV_X1    g295(.A(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n486_), .A2(new_n433_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n431_), .A3(new_n493_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n426_), .B(new_n501_), .C1(new_n420_), .C2(new_n419_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n495_), .A2(KEYINPUT95), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT95), .B1(new_n495_), .B2(new_n503_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT93), .B1(new_n412_), .B2(new_n417_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n398_), .A2(new_n402_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n409_), .A2(new_n411_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n417_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n431_), .B1(new_n499_), .B2(new_n493_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT33), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n509_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n418_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n490_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT96), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n492_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n497_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n492_), .A2(new_n518_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n431_), .B(new_n517_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n511_), .A2(new_n513_), .A3(new_n516_), .A4(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n502_), .B1(new_n506_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G22gat), .B(G50gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT28), .Z(new_n526_));
  NOR2_X1   g325(.A1(new_n484_), .A2(new_n485_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n528_), .A3(new_n526_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT88), .B1(new_n534_), .B2(new_n529_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G228gat), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n348_), .B1(KEYINPUT87), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT29), .B1(new_n484_), .B2(new_n485_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G78gat), .ZN(new_n541_));
  INV_X1    g340(.A(G78gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n542_), .A3(new_n539_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n537_), .A2(KEYINPUT87), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n210_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n546_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n533_), .B(new_n535_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n533_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n547_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G71gat), .B(G99gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G227gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G15gat), .B(G43gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n370_), .A2(KEYINPUT30), .A3(new_n380_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT30), .B1(new_n370_), .B2(new_n380_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n560_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n559_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n483_), .B(KEYINPUT31), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(KEYINPUT81), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n567_), .A3(new_n559_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n570_), .B(KEYINPUT81), .Z(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(new_n568_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n555_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n491_), .A2(new_n494_), .A3(new_n432_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n512_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n495_), .A2(new_n500_), .A3(KEYINPUT98), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n425_), .A2(new_n418_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n585_), .A2(KEYINPUT27), .A3(new_n510_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n516_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT27), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n535_), .A2(new_n533_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n551_), .B2(new_n547_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n548_), .A2(new_n549_), .A3(new_n533_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n573_), .B(new_n576_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n577_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n524_), .A2(new_n579_), .B1(new_n590_), .B2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n338_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT37), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(KEYINPUT72), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n245_), .A2(new_n322_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n235_), .A2(new_n244_), .A3(new_n295_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT35), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT70), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n235_), .A2(new_n295_), .A3(new_n244_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n235_), .A2(new_n244_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT34), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT34), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n615_), .B(new_n621_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n619_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n614_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n620_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n621_), .B1(new_n611_), .B2(new_n615_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n622_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n619_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(KEYINPUT35), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n608_), .B1(new_n625_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT71), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n625_), .B2(new_n631_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n635_), .ZN(new_n637_));
  AOI221_X4 g436(.A(new_n633_), .B1(new_n637_), .B2(new_n608_), .C1(new_n625_), .C2(new_n631_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n601_), .B(new_n604_), .C1(new_n636_), .C2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n608_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n623_), .A2(new_n624_), .A3(new_n612_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n613_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT71), .B1(new_n641_), .B2(new_n642_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n637_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n634_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(KEYINPUT72), .A4(new_n602_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n639_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n311_), .ZN(new_n649_));
  INV_X1    g448(.A(G231gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(new_n267_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n311_), .A2(G231gat), .A3(G233gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n258_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n259_), .A3(new_n652_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT74), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G127gat), .B(G155gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT16), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(new_n351_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(G211gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT17), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n658_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n658_), .A2(new_n664_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n656_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n663_), .A2(KEYINPUT17), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n665_), .A2(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n648_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n598_), .A2(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(G1gat), .A3(new_n584_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(KEYINPUT38), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(KEYINPUT38), .ZN(new_n674_));
  INV_X1    g473(.A(G1gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n645_), .A2(new_n646_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n597_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n669_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n337_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n584_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n673_), .B(new_n674_), .C1(new_n675_), .C2(new_n681_), .ZN(G1324gat));
  INV_X1    g481(.A(new_n589_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT99), .B1(new_n679_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(G8gat), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT39), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n679_), .A2(KEYINPUT99), .A3(new_n683_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n683_), .A2(new_n685_), .ZN(new_n691_));
  OAI22_X1  g490(.A1(new_n689_), .A2(new_n690_), .B1(new_n671_), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g492(.A1(new_n679_), .A2(new_n578_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G15gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n671_), .A2(G15gat), .A3(new_n577_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(G1326gat));
  XNOR2_X1  g499(.A(new_n554_), .B(KEYINPUT101), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n679_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G22gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT42), .ZN(new_n704_));
  INV_X1    g503(.A(new_n701_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(G22gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n671_), .B2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT102), .Z(G1327gat));
  NAND2_X1  g507(.A1(new_n524_), .A2(new_n579_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n590_), .A2(new_n596_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n669_), .A3(new_n676_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n338_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n680_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT69), .B1(new_n285_), .B2(new_n281_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n282_), .A2(new_n202_), .A3(new_n283_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n669_), .B(new_n335_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n287_), .A2(KEYINPUT103), .A3(new_n669_), .A4(new_n335_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n600_), .B(new_n603_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n723_));
  AND4_X1   g522(.A1(KEYINPUT72), .A2(new_n645_), .A3(new_n646_), .A4(new_n602_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n711_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT43), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n648_), .A2(new_n727_), .A3(new_n711_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n722_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n730_));
  OAI21_X1  g529(.A(new_n715_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n720_), .A2(new_n721_), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT43), .B(new_n597_), .C1(new_n647_), .C2(new_n639_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n727_), .B1(new_n648_), .B2(new_n711_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n730_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT105), .A3(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n731_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT44), .B(new_n732_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n740_), .A2(G29gat), .A3(new_n680_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n714_), .B1(new_n739_), .B2(new_n741_), .ZN(G1328gat));
  NOR4_X1   g541(.A1(new_n338_), .A2(new_n712_), .A3(G36gat), .A4(new_n589_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT108), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n743_), .B(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n740_), .A2(new_n683_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n731_), .B2(new_n737_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n749_));
  OAI21_X1  g548(.A(G36gat), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT106), .B(new_n747_), .C1(new_n731_), .C2(new_n737_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT46), .B(new_n746_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1329gat));
  NAND3_X1  g555(.A1(new_n740_), .A2(G43gat), .A3(new_n578_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n338_), .A2(new_n712_), .A3(new_n577_), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n738_), .A2(new_n757_), .B1(G43gat), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n713_), .B2(new_n701_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n740_), .A2(G50gat), .A3(new_n555_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n739_), .B2(new_n762_), .ZN(G1331gat));
  NOR2_X1   g562(.A1(new_n287_), .A2(new_n335_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(new_n669_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n677_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n584_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n765_), .A2(new_n597_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n670_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n680_), .A2(new_n249_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(G1332gat));
  INV_X1    g571(.A(new_n770_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(new_n251_), .A3(new_n683_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G64gat), .B1(new_n767_), .B2(new_n589_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n775_), .A2(KEYINPUT109), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(KEYINPUT109), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(KEYINPUT48), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT48), .B1(new_n776_), .B2(new_n777_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n774_), .B1(new_n778_), .B2(new_n779_), .ZN(G1333gat));
  OR3_X1    g579(.A1(new_n770_), .A2(G71gat), .A3(new_n577_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G71gat), .B1(new_n767_), .B2(new_n577_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n782_), .A2(new_n783_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1334gat));
  OAI21_X1  g585(.A(G78gat), .B1(new_n767_), .B2(new_n705_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT50), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n773_), .A2(new_n542_), .A3(new_n701_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1335gat));
  NOR2_X1   g589(.A1(new_n712_), .A2(new_n765_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n680_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT111), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n678_), .B(new_n765_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n584_), .A2(new_n213_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT112), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n794_), .B2(new_n796_), .ZN(G1336gat));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n214_), .A3(new_n683_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n794_), .A2(new_n683_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n214_), .ZN(G1337gat));
  AOI21_X1  g599(.A(new_n237_), .B1(new_n794_), .B2(new_n578_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n578_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n791_), .B2(new_n802_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g603(.A1(new_n791_), .A2(new_n210_), .A3(new_n555_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n765_), .A2(new_n678_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n555_), .B(new_n806_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G106gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT113), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n811_), .A3(G106gat), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n809_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n810_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n805_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT53), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n817_), .B(new_n805_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1339gat));
  NOR3_X1   g618(.A1(new_n335_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n639_), .A2(new_n678_), .A3(new_n647_), .A4(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n723_), .A2(new_n724_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n314_), .A2(new_n315_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n323_), .A2(new_n312_), .A3(new_n316_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n333_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n206_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n271_), .A2(new_n277_), .A3(new_n828_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n331_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n245_), .A2(new_n259_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n208_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n262_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n245_), .A2(new_n259_), .A3(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n833_), .A2(new_n270_), .A3(KEYINPUT55), .A4(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n264_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n270_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n276_), .B2(new_n208_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n265_), .A2(new_n269_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n268_), .B1(new_n841_), .B2(new_n275_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n838_), .A2(new_n839_), .A3(new_n843_), .A4(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(KEYINPUT56), .A3(new_n206_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n845_), .B2(new_n206_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  AOI211_X1 g648(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n845_), .C2(new_n206_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n830_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n824_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n331_), .A2(new_n827_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(KEYINPUT117), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n845_), .B2(new_n206_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n860_), .A2(new_n862_), .B1(new_n846_), .B2(KEYINPUT117), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n845_), .A2(new_n206_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n859_), .B1(new_n864_), .B2(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n335_), .A2(new_n829_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n857_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n855_), .B1(new_n869_), .B2(new_n676_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n676_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n865_), .B2(new_n863_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n871_), .B(KEYINPUT57), .C1(new_n872_), .C2(new_n857_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n669_), .B1(new_n854_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n823_), .B1(new_n875_), .B2(KEYINPUT120), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(KEYINPUT120), .B2(new_n875_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n683_), .A2(new_n594_), .A3(new_n584_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n823_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n851_), .B(KEYINPUT58), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n882_), .A2(new_n648_), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n882_), .B2(new_n648_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n874_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n881_), .B1(new_n886_), .B2(new_n678_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n879_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n880_), .B1(new_n878_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G113gat), .B1(new_n890_), .B2(new_n336_), .ZN(new_n891_));
  OR3_X1    g690(.A1(new_n888_), .A2(G113gat), .A3(new_n336_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1340gat));
  OAI21_X1  g692(.A(G120gat), .B1(new_n890_), .B2(new_n287_), .ZN(new_n894_));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n287_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n889_), .B(new_n896_), .C1(KEYINPUT60), .C2(new_n895_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(G1341gat));
  OAI21_X1  g697(.A(G127gat), .B1(new_n890_), .B2(new_n669_), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n888_), .A2(G127gat), .A3(new_n669_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1342gat));
  OAI21_X1  g700(.A(G134gat), .B1(new_n890_), .B2(new_n824_), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n888_), .A2(G134gat), .A3(new_n871_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1343gat));
  NOR3_X1   g703(.A1(new_n683_), .A2(new_n595_), .A3(new_n584_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT121), .Z(new_n906_));
  NAND2_X1  g705(.A1(new_n887_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n335_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n288_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g711(.A1(new_n907_), .A2(new_n669_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT61), .B(G155gat), .Z(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n908_), .B2(new_n676_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n648_), .A2(G162gat), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT122), .Z(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n908_), .B2(new_n918_), .ZN(G1347gat));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n680_), .A2(new_n577_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n683_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n701_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n877_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n336_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n920_), .B1(new_n925_), .B2(new_n362_), .ZN(new_n926_));
  OAI211_X1 g725(.A(KEYINPUT62), .B(G169gat), .C1(new_n924_), .C2(new_n336_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(G1348gat));
  INV_X1    g728(.A(new_n924_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G176gat), .B1(new_n930_), .B2(new_n288_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT119), .B1(new_n824_), .B2(new_n853_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n870_), .A2(new_n873_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n882_), .A2(new_n648_), .A3(new_n883_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n823_), .B1(new_n935_), .B2(new_n669_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n555_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n922_), .A2(new_n287_), .A3(new_n366_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n931_), .B1(new_n937_), .B2(new_n938_), .ZN(G1349gat));
  NOR3_X1   g738(.A1(new_n924_), .A2(new_n669_), .A3(new_n372_), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n937_), .A2(new_n678_), .A3(new_n683_), .A4(new_n921_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n941_), .A2(KEYINPUT123), .ZN(new_n942_));
  AOI21_X1  g741(.A(G183gat), .B1(new_n941_), .B2(KEYINPUT123), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n924_), .B2(new_n824_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n676_), .A2(new_n385_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n924_), .B2(new_n946_), .ZN(G1351gat));
  OR3_X1    g746(.A1(new_n680_), .A2(KEYINPUT124), .A3(new_n595_), .ZN(new_n948_));
  OAI21_X1  g747(.A(KEYINPUT124), .B1(new_n680_), .B2(new_n595_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n948_), .A2(new_n683_), .A3(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(KEYINPUT125), .B1(new_n887_), .B2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n936_), .A2(new_n953_), .A3(new_n950_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n335_), .B1(new_n952_), .B2(new_n954_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n955_), .A2(KEYINPUT126), .A3(new_n327_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n953_), .B1(new_n936_), .B2(new_n950_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n885_), .A2(new_n874_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n678_), .B1(new_n958_), .B2(new_n934_), .ZN(new_n959_));
  OAI211_X1 g758(.A(KEYINPUT125), .B(new_n951_), .C1(new_n959_), .C2(new_n823_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n336_), .B1(new_n957_), .B2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(G197gat), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n963_), .B1(new_n961_), .B2(G197gat), .ZN(new_n964_));
  AND3_X1   g763(.A1(new_n956_), .A2(new_n962_), .A3(new_n964_), .ZN(G1352gat));
  NAND2_X1  g764(.A1(new_n957_), .A2(new_n960_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n288_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g767(.A(new_n669_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n966_), .A2(new_n969_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(KEYINPUT127), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n970_), .B(new_n972_), .ZN(G1354gat));
  INV_X1    g772(.A(new_n966_), .ZN(new_n974_));
  OAI21_X1  g773(.A(G218gat), .B1(new_n974_), .B2(new_n824_), .ZN(new_n975_));
  INV_X1    g774(.A(G218gat), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n966_), .A2(new_n976_), .A3(new_n676_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n977_), .ZN(G1355gat));
endmodule


