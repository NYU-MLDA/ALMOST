//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT25), .B(G183gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT93), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT23), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n206_), .A2(new_n221_), .A3(new_n211_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n213_), .A2(new_n219_), .A3(new_n220_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT83), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n224_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n216_), .A3(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(G183gat), .B2(G190gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT22), .B(G169gat), .Z(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(G176gat), .B2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n210_), .B(KEYINPUT94), .Z(new_n231_));
  OAI21_X1  g030(.A(new_n223_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G197gat), .B(G204gat), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT21), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(new_n233_), .B2(KEYINPUT21), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n235_), .B(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n203_), .B1(new_n232_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G226gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT19), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n219_), .B1(G183gat), .B2(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT22), .B1(new_n207_), .B2(KEYINPUT84), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n208_), .B(new_n244_), .C1(new_n245_), .C2(KEYINPUT84), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n210_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n206_), .A2(KEYINPUT82), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n227_), .A2(new_n248_), .A3(new_n211_), .A4(new_n220_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n206_), .A2(KEYINPUT82), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n247_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT85), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(new_n247_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n237_), .B(new_n234_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n239_), .A2(new_n242_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT20), .B1(new_n232_), .B2(new_n238_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n254_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n238_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n257_), .B1(new_n260_), .B2(new_n242_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G8gat), .B(G36gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT96), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n202_), .B1(new_n261_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n258_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n259_), .A2(new_n238_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n241_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n239_), .A2(new_n241_), .A3(new_n256_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n267_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT100), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n260_), .B2(new_n241_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT100), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n267_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n269_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n268_), .B(new_n273_), .C1(new_n260_), .C2(new_n241_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n202_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT3), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT2), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n286_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n291_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n290_), .A2(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G22gat), .B(G50gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT28), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n299_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G78gat), .B(G106gat), .Z(new_n304_));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n238_), .B(new_n305_), .C1(new_n298_), .C2(new_n297_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n290_), .A2(new_n293_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n295_), .A2(new_n296_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n298_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT90), .B1(new_n309_), .B2(new_n255_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G228gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(G228gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(G233gat), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n306_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n306_), .B2(new_n310_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n304_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n317_), .A2(new_n318_), .A3(new_n304_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT91), .B(new_n304_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n324_));
  AND4_X1   g123(.A1(new_n303_), .A2(new_n321_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n319_), .B1(new_n322_), .B2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(KEYINPUT92), .B(new_n304_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n303_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n285_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT87), .B(G127gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G134gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(G113gat), .B(G120gat), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G134gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n332_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n339_), .A3(KEYINPUT31), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT31), .B1(new_n335_), .B2(new_n339_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT86), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT86), .B(new_n344_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n259_), .A2(KEYINPUT30), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n259_), .A2(KEYINPUT30), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n346_), .B(new_n347_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n347_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n348_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G71gat), .B(G99gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G15gat), .B(G43gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n335_), .A2(new_n339_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n307_), .A2(new_n308_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n297_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT97), .B1(new_n364_), .B2(KEYINPUT4), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT97), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n362_), .A2(new_n369_), .A3(new_n370_), .A4(new_n363_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n367_), .B1(new_n373_), .B2(new_n365_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G1gat), .B(G29gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(G57gat), .B(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n367_), .B(new_n379_), .C1(new_n373_), .C2(new_n365_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n361_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n331_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n359_), .A2(new_n360_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n351_), .A2(new_n354_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n357_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT88), .B1(new_n390_), .B2(new_n358_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n383_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n330_), .A2(new_n280_), .A3(new_n393_), .A4(new_n283_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n277_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n395_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n261_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n398_), .A3(new_n383_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n368_), .A2(new_n372_), .A3(new_n365_), .A4(new_n371_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n364_), .A2(new_n366_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n401_), .B(new_n380_), .C1(new_n365_), .C2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n275_), .A2(new_n281_), .A3(new_n400_), .A4(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n382_), .B(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n399_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n329_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n321_), .A2(new_n323_), .A3(new_n303_), .A4(new_n324_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  AOI211_X1 g210(.A(KEYINPUT101), .B(new_n392_), .C1(new_n394_), .C2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT101), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n394_), .A2(new_n411_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n392_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n385_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT64), .ZN(new_n418_));
  INV_X1    g217(.A(G99gat), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(KEYINPUT10), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(KEYINPUT10), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n418_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT10), .B(G99gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT64), .ZN(new_n424_));
  AOI21_X1  g223(.A(G106gat), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT66), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT6), .ZN(new_n429_));
  AND2_X1   g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G85gat), .A2(G92gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT9), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n434_), .A2(KEYINPUT65), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n434_), .B2(KEYINPUT65), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G85gat), .A2(G92gat), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n425_), .A2(new_n433_), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G85gat), .B(G92gat), .Z(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT68), .B(KEYINPUT8), .Z(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT67), .B(new_n444_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n430_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n453_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n430_), .A3(new_n454_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n444_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n448_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT8), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n440_), .B1(new_n452_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G29gat), .B(G36gat), .ZN(new_n464_));
  INV_X1    g263(.A(G43gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G50gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n464_), .B(G43gat), .ZN(new_n468_));
  INV_X1    g267(.A(G50gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G232gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT34), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n463_), .A2(new_n471_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n467_), .A2(new_n470_), .A3(KEYINPUT15), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT15), .B1(new_n467_), .B2(new_n470_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(new_n463_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n475_), .A2(new_n472_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n477_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G190gat), .B(G218gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G134gat), .ZN(new_n486_));
  INV_X1    g285(.A(G162gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT76), .Z(new_n491_));
  OR2_X1    g290(.A1(new_n478_), .A2(new_n479_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n463_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(KEYINPUT74), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT74), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n480_), .B2(new_n463_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n476_), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(KEYINPUT75), .A3(new_n482_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT75), .B1(new_n497_), .B2(new_n482_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n484_), .B(new_n491_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT37), .ZN(new_n502_));
  INV_X1    g301(.A(new_n500_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n483_), .B1(new_n503_), .B2(new_n498_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n488_), .B(KEYINPUT36), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n501_), .B(new_n502_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n484_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n505_), .B(KEYINPUT77), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n502_), .B1(new_n511_), .B2(new_n501_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G127gat), .B(G155gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G183gat), .B(G211gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G71gat), .B(G78gat), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n522_), .A3(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G231gat), .A2(G233gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT78), .ZN(new_n529_));
  INV_X1    g328(.A(G1gat), .ZN(new_n530_));
  INV_X1    g329(.A(G8gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G1gat), .B(G8gat), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n529_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n527_), .B(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n518_), .B1(new_n542_), .B2(KEYINPUT80), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n542_), .B2(new_n518_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(new_n543_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n513_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n463_), .A2(new_n525_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n463_), .A2(new_n525_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G120gat), .B(G148gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n463_), .B2(new_n525_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT12), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n561_), .B(new_n564_), .C1(new_n463_), .C2(new_n525_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n563_), .A2(new_n552_), .A3(new_n550_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n554_), .B(new_n560_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n563_), .A2(new_n565_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n571_), .A2(KEYINPUT71), .A3(new_n550_), .A4(new_n552_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n567_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n553_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n559_), .B(KEYINPUT73), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n570_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT13), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n471_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n467_), .A2(new_n470_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n541_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n585_), .A3(KEYINPUT81), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT81), .B1(new_n583_), .B2(new_n585_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n582_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n492_), .A2(new_n541_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n583_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n582_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G113gat), .B(G141gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n207_), .ZN(new_n594_));
  INV_X1    g393(.A(G197gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n589_), .B(new_n598_), .C1(new_n591_), .C2(new_n582_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n580_), .A2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n417_), .A2(new_n549_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n530_), .A3(new_n383_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT102), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n501_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n548_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n417_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n602_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n393_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n607_), .B(new_n612_), .C1(new_n605_), .C2(new_n604_), .ZN(G1324gat));
  AND2_X1   g412(.A1(new_n610_), .A2(new_n602_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n285_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G8gat), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(KEYINPUT103), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(KEYINPUT103), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n617_), .A2(KEYINPUT103), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n615_), .A2(G8gat), .A3(new_n619_), .A4(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n603_), .A2(new_n531_), .A3(new_n285_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n618_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1325gat));
  INV_X1    g424(.A(G15gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n614_), .B2(new_n392_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT41), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n603_), .A2(new_n626_), .A3(new_n392_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1326gat));
  INV_X1    g429(.A(G22gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n603_), .A2(new_n631_), .A3(new_n330_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G22gat), .B1(new_n611_), .B2(new_n410_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(KEYINPUT42), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT42), .B1(new_n634_), .B2(new_n635_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n632_), .B1(new_n636_), .B2(new_n637_), .ZN(G1327gat));
  NOR3_X1   g437(.A1(new_n580_), .A2(new_n609_), .A3(new_n601_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n417_), .A2(new_n640_), .A3(new_n513_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n417_), .B2(new_n513_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n639_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n414_), .A2(new_n415_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT101), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n414_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n647_), .A2(new_n648_), .B1(new_n331_), .B2(new_n384_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n513_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT43), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n417_), .A2(new_n640_), .A3(new_n513_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n644_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n639_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n645_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n393_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n649_), .A2(new_n608_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(new_n639_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(G29gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n393_), .B2(new_n661_), .ZN(G1328gat));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n663_), .A3(new_n285_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT45), .ZN(new_n665_));
  OAI21_X1  g464(.A(G36gat), .B1(new_n656_), .B2(new_n284_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1329gat));
  OAI21_X1  g468(.A(new_n465_), .B1(new_n660_), .B2(new_n415_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n361_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G43gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n656_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g473(.A(G50gat), .B1(new_n656_), .B2(new_n410_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n659_), .A2(new_n469_), .A3(new_n330_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1331gat));
  NAND3_X1  g476(.A1(new_n610_), .A2(new_n601_), .A3(new_n580_), .ZN(new_n678_));
  INV_X1    g477(.A(G57gat), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n393_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n579_), .A2(new_n513_), .A3(new_n548_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n600_), .B(new_n649_), .C1(KEYINPUT106), .C2(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(KEYINPUT106), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n393_), .B1(new_n685_), .B2(KEYINPUT107), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(KEYINPUT107), .B2(new_n685_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n680_), .B1(new_n687_), .B2(new_n679_), .ZN(G1332gat));
  OAI21_X1  g487(.A(G64gat), .B1(new_n678_), .B2(new_n284_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT48), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n284_), .A2(G64gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n684_), .B2(new_n691_), .ZN(G1333gat));
  OAI21_X1  g491(.A(G71gat), .B1(new_n678_), .B2(new_n415_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT49), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n684_), .A2(G71gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n415_), .B2(new_n695_), .ZN(G1334gat));
  OAI21_X1  g495(.A(G78gat), .B1(new_n678_), .B2(new_n410_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT50), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n684_), .A2(G78gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n410_), .B2(new_n699_), .ZN(G1335gat));
  NOR3_X1   g499(.A1(new_n579_), .A2(new_n609_), .A3(new_n600_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n658_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n383_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT108), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n653_), .A2(new_n701_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n383_), .A2(G85gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(G1336gat));
  AOI21_X1  g507(.A(G92gat), .B1(new_n703_), .B2(new_n285_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n285_), .A2(G92gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n706_), .B2(new_n710_), .ZN(G1337gat));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n392_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n361_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n712_), .A2(G99gat), .B1(new_n703_), .B2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n330_), .B(new_n701_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT109), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n653_), .A2(new_n719_), .A3(new_n330_), .A4(new_n701_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n720_), .A3(G106gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT52), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n718_), .A2(new_n720_), .A3(new_n723_), .A4(G106gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n702_), .A2(G106gat), .A3(new_n410_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n716_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n716_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n729_), .B(new_n726_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1339gat));
  NAND3_X1  g530(.A1(new_n549_), .A2(new_n601_), .A3(new_n579_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT54), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n736_), .B2(new_n732_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n600_), .A2(new_n570_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n563_), .A2(new_n552_), .A3(new_n565_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n550_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(new_n741_), .B2(new_n566_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n742_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n575_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT56), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n751_), .B(new_n575_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n740_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n583_), .A2(new_n585_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT81), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n582_), .B1(new_n757_), .B2(new_n586_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n758_), .B2(new_n598_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n581_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(KEYINPUT112), .A3(new_n596_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n590_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(new_n599_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n572_), .A2(new_n573_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n575_), .B1(new_n765_), .B2(new_n554_), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n553_), .B(new_n559_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n576_), .A2(KEYINPUT113), .A3(new_n764_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n753_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n772_), .A2(KEYINPUT57), .A3(new_n608_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT57), .B1(new_n772_), .B2(new_n608_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n738_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n764_), .A2(new_n570_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT55), .B1(new_n572_), .B2(new_n573_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n749_), .B1(new_n777_), .B2(new_n746_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n751_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n748_), .A2(KEYINPUT56), .A3(new_n749_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n513_), .B1(new_n781_), .B2(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(KEYINPUT58), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n513_), .B(new_n785_), .C1(new_n781_), .C2(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n784_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n770_), .A2(new_n771_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n739_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n608_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n738_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n775_), .A2(new_n787_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n737_), .B1(new_n794_), .B2(new_n548_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n331_), .A2(new_n383_), .A3(new_n671_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT59), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(KEYINPUT59), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n791_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n772_), .A2(KEYINPUT57), .A3(new_n608_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n609_), .B1(new_n802_), .B2(new_n787_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n798_), .B1(new_n803_), .B2(new_n737_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n797_), .A2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT118), .B(G113gat), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n601_), .A2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT119), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n796_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n792_), .B1(new_n801_), .B2(new_n738_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n609_), .B1(new_n813_), .B2(new_n787_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT116), .B(new_n812_), .C1(new_n814_), .C2(new_n737_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n600_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n601_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT117), .B1(new_n821_), .B2(G113gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n809_), .B1(new_n820_), .B2(new_n822_), .ZN(G1340gat));
  OAI21_X1  g622(.A(G120gat), .B1(new_n805_), .B2(new_n579_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n579_), .B2(KEYINPUT60), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(KEYINPUT60), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AND4_X1   g628(.A1(new_n825_), .A2(new_n816_), .A3(new_n827_), .A4(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n825_), .B1(new_n831_), .B2(new_n827_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n824_), .B1(new_n830_), .B2(new_n832_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n816_), .B2(new_n609_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n797_), .A2(G127gat), .A3(new_n804_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n609_), .ZN(G1342gat));
  NOR3_X1   g635(.A1(new_n805_), .A2(new_n336_), .A3(new_n650_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n608_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n816_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT121), .A3(new_n336_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n608_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(G134gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n837_), .B1(new_n840_), .B2(new_n843_), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n795_), .A2(new_n393_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n285_), .A2(new_n392_), .A3(new_n410_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n601_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT122), .B(G141gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT123), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n848_), .B(new_n850_), .ZN(G1344gat));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n580_), .A3(new_n846_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g652(.A1(new_n847_), .A2(new_n548_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT61), .B(G155gat), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  NAND4_X1  g655(.A1(new_n845_), .A2(G162gat), .A3(new_n513_), .A4(new_n846_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n794_), .A2(new_n548_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n737_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AND4_X1   g659(.A1(new_n383_), .A2(new_n860_), .A3(new_n838_), .A4(new_n846_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n857_), .B1(new_n861_), .B2(G162gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT124), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n857_), .B(new_n864_), .C1(new_n861_), .C2(G162gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n284_), .A2(new_n383_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n415_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n410_), .B(new_n869_), .C1(new_n803_), .C2(new_n737_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870_), .B2(new_n601_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT125), .B(G169gat), .C1(new_n870_), .C2(new_n601_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(KEYINPUT62), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n871_), .A2(new_n872_), .A3(new_n876_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n870_), .A2(new_n601_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n875_), .B(new_n877_), .C1(new_n229_), .C2(new_n878_), .ZN(G1348gat));
  NOR2_X1   g678(.A1(new_n795_), .A2(new_n330_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n880_), .A2(G176gat), .A3(new_n580_), .A4(new_n869_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n208_), .B1(new_n870_), .B2(new_n579_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(KEYINPUT126), .A3(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1349gat));
  NOR3_X1   g686(.A1(new_n870_), .A2(new_n548_), .A3(new_n204_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n880_), .A2(new_n609_), .A3(new_n869_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n214_), .ZN(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n870_), .B2(new_n650_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n838_), .A2(new_n205_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n870_), .B2(new_n892_), .ZN(G1351gat));
  NOR4_X1   g692(.A1(new_n795_), .A2(new_n392_), .A3(new_n410_), .A4(new_n868_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n600_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g695(.A1(new_n860_), .A2(new_n415_), .A3(new_n330_), .A4(new_n867_), .ZN(new_n897_));
  OAI22_X1  g696(.A1(new_n897_), .A2(new_n579_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n897_), .A2(new_n579_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1353gat));
  AOI211_X1 g701(.A(KEYINPUT63), .B(G211gat), .C1(new_n894_), .C2(new_n609_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT63), .B(G211gat), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n897_), .A2(new_n548_), .A3(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1354gat));
  AND3_X1   g705(.A1(new_n894_), .A2(G218gat), .A3(new_n513_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G218gat), .B1(new_n894_), .B2(new_n838_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1355gat));
endmodule


