//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203_));
  INV_X1    g002(.A(G85gat), .ZN(new_n204_));
  INV_X1    g003(.A(G92gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n203_), .B(new_n206_), .C1(new_n208_), .C2(KEYINPUT64), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n206_), .A2(new_n210_), .A3(KEYINPUT9), .A4(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n209_), .A2(new_n211_), .A3(new_n216_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n206_), .A2(new_n207_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI211_X1 g025(.A(KEYINPUT8), .B(new_n222_), .C1(new_n226_), .C2(new_n216_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  INV_X1    g028(.A(G99gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n218_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n223_), .B(new_n231_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n222_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n228_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n221_), .B1(new_n227_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(new_n221_), .C1(new_n227_), .C2(new_n236_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  INV_X1    g040(.A(G78gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G71gat), .ZN(new_n243_));
  INV_X1    g042(.A(G71gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G78gat), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n241_), .A2(KEYINPUT11), .A3(new_n243_), .A4(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G64gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G57gat), .ZN(new_n248_));
  INV_X1    g047(.A(G57gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G64gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n250_), .A3(KEYINPUT11), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n243_), .A2(new_n245_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n254_));
  OAI211_X1 g053(.A(KEYINPUT67), .B(new_n246_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT12), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n248_), .A2(new_n250_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT67), .B1(new_n260_), .B2(new_n246_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n238_), .A2(new_n240_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n246_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n237_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT12), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n221_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n234_), .A2(new_n235_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT8), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n234_), .A2(new_n228_), .A3(new_n235_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n270_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n269_), .B1(new_n274_), .B2(new_n264_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n263_), .A2(new_n268_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n263_), .A2(new_n268_), .A3(KEYINPUT68), .A4(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n264_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n266_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n282_), .B(new_n269_), .C1(new_n281_), .C2(new_n266_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n279_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT5), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT69), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n278_), .A2(new_n283_), .A3(new_n279_), .A4(new_n288_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n291_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n298_), .B(new_n291_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n297_), .A2(KEYINPUT13), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT13), .B1(new_n297_), .B2(new_n299_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n202_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT13), .ZN(new_n303_));
  INV_X1    g102(.A(new_n299_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n292_), .B(new_n293_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n298_), .B1(new_n305_), .B2(new_n291_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n303_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n297_), .A2(KEYINPUT13), .A3(new_n299_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT72), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G29gat), .B(G36gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G43gat), .B(G50gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT15), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n238_), .A2(new_n315_), .A3(new_n240_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT35), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G232gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT34), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n274_), .A2(new_n314_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n320_), .A2(new_n317_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G190gat), .B(G218gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G134gat), .B(G162gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  OR4_X1    g127(.A1(KEYINPUT36), .A2(new_n324_), .A3(new_n325_), .A4(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n328_), .B(KEYINPUT36), .Z(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT37), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT37), .A4(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G15gat), .B(G22gat), .ZN(new_n338_));
  INV_X1    g137(.A(G1gat), .ZN(new_n339_));
  INV_X1    g138(.A(G8gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT14), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G8gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G231gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n265_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n344_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(new_n345_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(G231gat), .B2(G233gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n264_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G155gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT16), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G183gat), .B(G211gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT17), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n352_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT74), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n359_), .A4(new_n353_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n359_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n357_), .A2(new_n358_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n367_), .A2(new_n347_), .A3(new_n351_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n337_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n311_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT99), .ZN(new_n375_));
  INV_X1    g174(.A(G134gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G127gat), .ZN(new_n377_));
  INV_X1    g176(.A(G127gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G134gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT83), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(KEYINPUT85), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(KEYINPUT85), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n383_), .A2(KEYINPUT83), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n377_), .A2(new_n379_), .A3(KEYINPUT83), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n385_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n382_), .A2(new_n384_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT84), .B1(new_n395_), .B2(new_n385_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n388_), .B(new_n389_), .C1(new_n394_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G141gat), .ZN(new_n398_));
  INV_X1    g197(.A(G148gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT86), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT1), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n403_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n404_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT1), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n406_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT87), .A3(new_n403_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n400_), .A2(KEYINPUT3), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT2), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n401_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n400_), .A2(KEYINPUT3), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n412_), .A2(new_n406_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n410_), .A2(new_n416_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n397_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT100), .B(KEYINPUT4), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT97), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n392_), .A2(new_n428_), .A3(new_n387_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n392_), .B2(new_n387_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT98), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n424_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n392_), .A2(new_n387_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT97), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n392_), .A2(new_n428_), .A3(new_n387_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n410_), .A2(new_n416_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n423_), .A2(new_n422_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT98), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n433_), .B1(new_n441_), .B2(new_n425_), .ZN(new_n442_));
  AOI211_X1 g241(.A(new_n375_), .B(new_n427_), .C1(KEYINPUT4), .C2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G85gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT0), .B(G57gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n442_), .B2(new_n375_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT101), .B1(new_n443_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n427_), .B1(new_n442_), .B2(KEYINPUT4), .ZN(new_n451_));
  INV_X1    g250(.A(new_n375_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT101), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n431_), .A2(new_n424_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(KEYINPUT98), .C1(new_n424_), .C2(new_n397_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n452_), .A3(new_n433_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n447_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT19), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n465_), .B(KEYINPUT93), .Z(new_n466_));
  NOR2_X1   g265(.A1(G169gat), .A2(G176gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT24), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G169gat), .A2(G176gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT24), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n471_), .B2(new_n467_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT26), .B(G190gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT95), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT25), .B(G183gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G183gat), .A2(G190gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT81), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(KEYINPUT77), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT77), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G183gat), .A3(G190gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n481_), .B1(new_n485_), .B2(new_n480_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(KEYINPUT81), .A4(KEYINPUT23), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n477_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT22), .B(G169gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT79), .B(G176gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n479_), .A2(new_n480_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n485_), .B2(new_n480_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G183gat), .A2(G190gat), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n470_), .B(new_n492_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT21), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT90), .B(G204gat), .ZN(new_n499_));
  INV_X1    g298(.A(G197gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G197gat), .A2(G204gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G211gat), .B(G218gat), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n500_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n498_), .B1(G197gat), .B2(G204gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n501_), .A2(new_n502_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n504_), .A2(KEYINPUT21), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n503_), .A2(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n497_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT22), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G169gat), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n514_), .A2(KEYINPUT78), .ZN(new_n515_));
  INV_X1    g314(.A(G169gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT22), .B1(new_n516_), .B2(KEYINPUT78), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n491_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT80), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT80), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n515_), .A2(new_n520_), .A3(new_n491_), .A4(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n486_), .B(new_n487_), .C1(G183gat), .C2(G190gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n470_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n494_), .A2(new_n472_), .ZN(new_n525_));
  INV_X1    g324(.A(G183gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT25), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(KEYINPUT25), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(KEYINPUT75), .B2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(KEYINPUT75), .ZN(new_n530_));
  INV_X1    g329(.A(G190gat), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n531_), .A2(KEYINPUT76), .A3(KEYINPUT26), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT26), .B1(new_n531_), .B2(KEYINPUT76), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n525_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT20), .B1(new_n536_), .B2(new_n511_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n512_), .B1(new_n537_), .B2(KEYINPUT94), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n519_), .A2(new_n521_), .B1(G169gat), .B2(G176gat), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n540_), .A2(new_n523_), .B1(new_n534_), .B2(new_n525_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n510_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n542_), .B2(KEYINPUT20), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n466_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n465_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n497_), .B2(new_n511_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n536_), .B2(new_n511_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n549_), .A3(KEYINPUT96), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT96), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT20), .B1(new_n541_), .B2(new_n510_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n546_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G8gat), .B(G36gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT18), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G64gat), .B(G92gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  AND3_X1   g357(.A1(new_n544_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n544_), .B2(new_n554_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n460_), .A2(KEYINPUT33), .A3(new_n447_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n456_), .A2(new_n463_), .A3(new_n561_), .A4(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT103), .ZN(new_n564_));
  INV_X1    g363(.A(new_n447_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n459_), .B(new_n565_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n461_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n460_), .A2(KEYINPUT103), .A3(new_n447_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n558_), .A2(KEYINPUT32), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n510_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n497_), .A2(KEYINPUT102), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n497_), .A2(KEYINPUT102), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n549_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n465_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n543_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n542_), .A2(new_n539_), .A3(KEYINPUT20), .ZN(new_n579_));
  INV_X1    g378(.A(new_n466_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .A4(new_n512_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n569_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n544_), .A2(new_n554_), .A3(new_n569_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n567_), .A2(new_n568_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n563_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n440_), .A2(KEYINPUT29), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n440_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(G228gat), .ZN(new_n592_));
  INV_X1    g391(.A(G233gat), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n510_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n594_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n440_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n571_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G78gat), .B(G106gat), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n440_), .B2(KEYINPUT29), .ZN(new_n606_));
  XOR2_X1   g405(.A(G22gat), .B(G50gat), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n609_));
  INV_X1    g408(.A(new_n605_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n424_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n606_), .A2(new_n608_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n608_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n511_), .A2(new_n597_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n602_), .B1(new_n616_), .B2(new_n600_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n604_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n604_), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G71gat), .B(G99gat), .ZN(new_n621_));
  INV_X1    g420(.A(G43gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT31), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G227gat), .A2(G233gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(G15gat), .Z(new_n629_));
  NOR2_X1   g428(.A1(new_n536_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n524_), .B2(new_n535_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n627_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n541_), .A2(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n536_), .A2(new_n629_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n626_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n633_), .A2(new_n636_), .A3(new_n397_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n397_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n625_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n397_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n630_), .A2(new_n632_), .A3(new_n627_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n626_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n633_), .A2(new_n636_), .A3(new_n397_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n624_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n620_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n586_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n614_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n603_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n616_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n604_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n639_), .A4(new_n645_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n637_), .A2(new_n638_), .A3(new_n625_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n624_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n618_), .A2(new_n619_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n654_), .A2(new_n657_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n561_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT27), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n559_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n558_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n577_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n581_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  AOI22_X1  g464(.A1(new_n659_), .A2(new_n660_), .B1(new_n661_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n648_), .A2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n344_), .B(new_n314_), .Z(new_n669_));
  NAND2_X1  g468(.A1(G229gat), .A2(G233gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n315_), .A2(new_n344_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n348_), .A2(new_n314_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n670_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(G113gat), .B(G141gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(G169gat), .B(G197gat), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n677_), .B(new_n678_), .Z(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n676_), .A2(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n668_), .A2(KEYINPUT104), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n586_), .A2(new_n647_), .B1(new_n658_), .B2(new_n666_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n684_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n685_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n567_), .A2(new_n568_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n373_), .A2(new_n690_), .A3(new_n339_), .A4(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT105), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT38), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n370_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n329_), .A2(new_n332_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n668_), .A2(new_n698_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n688_), .B1(new_n302_), .B2(new_n309_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G1gat), .B1(new_n704_), .B2(new_n691_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n696_), .A2(new_n697_), .A3(new_n705_), .ZN(G1324gat));
  INV_X1    g505(.A(new_n666_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n373_), .A2(new_n690_), .A3(new_n340_), .A4(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n707_), .A3(new_n703_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(G8gat), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G8gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g513(.A1(new_n702_), .A2(new_n646_), .A3(new_n703_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(G15gat), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n717_), .A2(new_n720_), .A3(new_n718_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n373_), .A2(new_n690_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n646_), .ZN(new_n725_));
  OR3_X1    g524(.A1(new_n724_), .A2(G15gat), .A3(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n723_), .A3(new_n726_), .ZN(G1326gat));
  INV_X1    g526(.A(new_n620_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G22gat), .B1(new_n704_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT42), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n728_), .A2(G22gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n724_), .B2(new_n731_), .ZN(G1327gat));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n703_), .A2(KEYINPUT109), .A3(new_n370_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n337_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT43), .B1(new_n687_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n737_));
  INV_X1    g536(.A(new_n667_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n647_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n563_), .B2(new_n585_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n737_), .B(new_n337_), .C1(new_n738_), .C2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n734_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT109), .B1(new_n703_), .B2(new_n370_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n733_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n703_), .A2(new_n370_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n748_), .A2(KEYINPUT44), .A3(new_n742_), .A4(new_n734_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n745_), .A2(G29gat), .A3(new_n692_), .A4(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(G29gat), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n700_), .A2(new_n698_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n302_), .B2(new_n309_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n690_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n755_), .B2(new_n691_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n750_), .A2(new_n756_), .ZN(G1328gat));
  NAND3_X1  g556(.A1(new_n745_), .A2(new_n707_), .A3(new_n749_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G36gat), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n666_), .A2(G36gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n690_), .A2(new_n754_), .A3(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n764_), .A3(KEYINPUT46), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(G36gat), .B2(new_n758_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT111), .B(KEYINPUT46), .Z(new_n767_));
  OAI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(G1329gat));
  NOR2_X1   g567(.A1(new_n725_), .A2(new_n622_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n745_), .A2(new_n749_), .A3(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n622_), .B1(new_n755_), .B2(new_n725_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g572(.A1(new_n755_), .A2(G50gat), .A3(new_n728_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n745_), .A2(new_n620_), .A3(new_n749_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n775_), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT112), .B1(new_n775_), .B2(G50gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(G1331gat));
  NOR2_X1   g577(.A1(new_n310_), .A2(new_n684_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n668_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(new_n372_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n249_), .A3(new_n692_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n702_), .A2(new_n779_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G57gat), .B1(new_n783_), .B2(new_n691_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1332gat));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n247_), .A3(new_n707_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n701_), .A2(new_n684_), .A3(new_n310_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n707_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n789_), .B2(G64gat), .ZN(new_n790_));
  AOI211_X1 g589(.A(KEYINPUT48), .B(new_n247_), .C1(new_n788_), .C2(new_n707_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n786_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1333gat));
  OAI21_X1  g593(.A(G71gat), .B1(new_n783_), .B2(new_n725_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT49), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n781_), .A2(new_n244_), .A3(new_n646_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1334gat));
  NAND3_X1  g597(.A1(new_n781_), .A2(new_n242_), .A3(new_n620_), .ZN(new_n799_));
  OAI21_X1  g598(.A(G78gat), .B1(new_n783_), .B2(new_n728_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(KEYINPUT50), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(KEYINPUT50), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n799_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT114), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n799_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1335gat));
  NOR2_X1   g606(.A1(new_n780_), .A2(new_n753_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n204_), .A3(new_n692_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n742_), .A2(new_n370_), .A3(new_n779_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n742_), .A2(new_n779_), .A3(KEYINPUT115), .A4(new_n370_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n691_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n809_), .B1(new_n814_), .B2(new_n204_), .ZN(G1336gat));
  NAND3_X1  g614(.A1(new_n808_), .A2(new_n205_), .A3(new_n707_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n666_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n205_), .ZN(G1337gat));
  AOI21_X1  g617(.A(new_n725_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n230_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n808_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n646_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT51), .B1(new_n820_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n825_));
  OAI221_X1 g624(.A(new_n825_), .B1(new_n821_), .B2(new_n822_), .C1(new_n819_), .C2(new_n230_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1338gat));
  NAND3_X1  g626(.A1(new_n808_), .A2(new_n218_), .A3(new_n620_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n742_), .A2(new_n779_), .A3(new_n620_), .A4(new_n370_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(G106gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n829_), .B2(G106gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n278_), .A2(new_n835_), .A3(new_n279_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n263_), .A2(new_n268_), .A3(new_n275_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n263_), .A2(new_n268_), .A3(new_n280_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n837_), .A2(KEYINPUT55), .B1(new_n838_), .B2(new_n269_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n290_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n842_), .B(new_n289_), .C1(new_n836_), .C2(new_n839_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n679_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(KEYINPUT118), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n670_), .B1(new_n348_), .B2(new_n314_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n673_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(KEYINPUT118), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n681_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT119), .B1(new_n844_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT58), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT119), .B(new_n854_), .C1(new_n844_), .C2(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n337_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n850_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n684_), .B(new_n305_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT57), .B(new_n700_), .C1(new_n858_), .C2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n850_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n699_), .B1(new_n862_), .B2(new_n859_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n856_), .B(new_n861_), .C1(new_n863_), .C2(KEYINPUT57), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT116), .B1(new_n370_), .B2(new_n684_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n688_), .A2(new_n866_), .A3(new_n366_), .A4(new_n369_), .ZN(new_n867_));
  AND4_X1   g666(.A1(new_n335_), .A2(new_n865_), .A3(new_n336_), .A4(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n868_), .A2(new_n307_), .A3(new_n308_), .A4(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n869_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n864_), .A2(new_n370_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n707_), .A2(new_n691_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n874_), .A2(new_n657_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877_), .B2(new_n684_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n856_), .A2(new_n861_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n862_), .A2(new_n859_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880_), .B2(new_n700_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n370_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n871_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n657_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n875_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(KEYINPUT59), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n884_), .A2(new_n885_), .A3(new_n875_), .A4(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n888_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n684_), .A2(G113gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT121), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n878_), .B1(new_n892_), .B2(new_n894_), .ZN(G1340gat));
  NAND3_X1  g694(.A1(new_n888_), .A2(new_n311_), .A3(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G120gat), .ZN(new_n897_));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n310_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(KEYINPUT60), .B2(new_n898_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n886_), .B2(new_n900_), .ZN(G1341gat));
  NOR4_X1   g700(.A1(new_n874_), .A2(new_n657_), .A3(new_n370_), .A4(new_n876_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT122), .B1(new_n902_), .B2(G127gat), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n370_), .A2(new_n378_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n887_), .A2(KEYINPUT59), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n891_), .B(new_n904_), .C1(new_n877_), .C2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(new_n378_), .C1(new_n886_), .C2(new_n370_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n903_), .A2(new_n906_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n903_), .A2(new_n906_), .A3(new_n908_), .A4(KEYINPUT123), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1342gat));
  OAI21_X1  g712(.A(new_n376_), .B1(new_n886_), .B2(new_n700_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n914_), .A2(KEYINPUT124), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n888_), .A2(G134gat), .A3(new_n337_), .A4(new_n891_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(KEYINPUT124), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(G1343gat));
  INV_X1    g717(.A(new_n654_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n884_), .A2(new_n919_), .A3(new_n875_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n688_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n398_), .ZN(G1344gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n310_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n399_), .ZN(G1345gat));
  NOR2_X1   g723(.A1(new_n920_), .A2(new_n370_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT61), .B(G155gat), .Z(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1346gat));
  INV_X1    g726(.A(G162gat), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n920_), .A2(new_n928_), .A3(new_n735_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n920_), .B2(new_n700_), .ZN(new_n930_));
  OR2_X1    g729(.A1(new_n930_), .A2(KEYINPUT125), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(KEYINPUT125), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n929_), .B1(new_n931_), .B2(new_n932_), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n666_), .A2(new_n692_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n934_), .A2(new_n885_), .A3(new_n684_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT126), .B1(new_n936_), .B2(new_n516_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n938_), .B(G169gat), .C1(new_n874_), .C2(new_n935_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n937_), .A2(KEYINPUT62), .A3(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941_));
  OAI211_X1 g740(.A(KEYINPUT126), .B(new_n941_), .C1(new_n936_), .C2(new_n516_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n936_), .A2(new_n490_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n940_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n940_), .A2(KEYINPUT127), .A3(new_n942_), .A4(new_n943_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1348gat));
  NAND2_X1  g747(.A1(new_n934_), .A2(new_n885_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n874_), .A2(new_n949_), .ZN(new_n950_));
  AND3_X1   g749(.A1(new_n950_), .A2(G176gat), .A3(new_n311_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n311_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n951_), .B1(new_n491_), .B2(new_n952_), .ZN(G1349gat));
  NAND2_X1  g752(.A1(new_n950_), .A2(new_n698_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n476_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n526_), .B2(new_n954_), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n950_), .A2(new_n475_), .A3(new_n699_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n874_), .A2(new_n735_), .A3(new_n949_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n531_), .ZN(G1351gat));
  AND3_X1   g758(.A1(new_n884_), .A2(new_n919_), .A3(new_n934_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n684_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n311_), .ZN(new_n963_));
  MUX2_X1   g762(.A(new_n499_), .B(G204gat), .S(new_n963_), .Z(G1353gat));
  NAND2_X1  g763(.A1(new_n960_), .A2(new_n698_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  AND2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n965_), .A2(new_n966_), .A3(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n968_), .B1(new_n965_), .B2(new_n966_), .ZN(G1354gat));
  INV_X1    g768(.A(G218gat), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n960_), .A2(new_n970_), .A3(new_n699_), .ZN(new_n971_));
  AND2_X1   g770(.A1(new_n960_), .A2(new_n337_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(new_n970_), .ZN(G1355gat));
endmodule


