//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT83), .ZN(new_n203_));
  INV_X1    g002(.A(G155gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n213_));
  INV_X1    g012(.A(G141gat), .ZN(new_n214_));
  INV_X1    g013(.A(G148gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n216_), .A2(new_n217_), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n206_), .A2(new_n207_), .B1(G155gat), .B2(G162gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n219_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT28), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n212_), .A2(new_n218_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G228gat), .A2(G233gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT87), .B(KEYINPUT21), .Z(new_n237_));
  INV_X1    g036(.A(KEYINPUT86), .ZN(new_n238_));
  INV_X1    g037(.A(G204gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(G197gat), .ZN(new_n240_));
  INV_X1    g039(.A(G197gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(G197gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT85), .ZN(new_n245_));
  OR3_X1    g044(.A1(new_n241_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n237_), .A2(new_n243_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(G204gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n244_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n248_), .A2(new_n250_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT84), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n235_), .A2(new_n236_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n236_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n264_));
  INV_X1    g063(.A(G78gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n258_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n233_), .B1(new_n219_), .B2(new_n228_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n247_), .A2(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n268_));
  OAI21_X1  g067(.A(G78gat), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(G106gat), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(G106gat), .B1(new_n266_), .B2(new_n269_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G22gat), .B(G50gat), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n266_), .A2(new_n269_), .ZN(new_n276_));
  INV_X1    g075(.A(G106gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n275_), .B1(new_n278_), .B2(new_n270_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n263_), .B1(new_n274_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n273_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n281_), .A2(new_n260_), .A3(new_n262_), .A4(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT25), .B(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT73), .B1(new_n285_), .B2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G190gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n284_), .B(new_n286_), .C1(new_n287_), .C2(KEYINPUT73), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT74), .ZN(new_n289_));
  INV_X1    g088(.A(G183gat), .ZN(new_n290_));
  INV_X1    g089(.A(G190gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT23), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n295_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n285_), .A2(G190gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n291_), .A2(KEYINPUT26), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n284_), .A4(new_n286_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n289_), .A2(new_n302_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G169gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT22), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G169gat), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G176gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT75), .A3(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n317_));
  OAI21_X1  g116(.A(G169gat), .B1(new_n317_), .B2(G176gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n292_), .A2(KEYINPUT76), .A3(new_n294_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n320_), .B(KEYINPUT23), .C1(new_n290_), .C2(new_n291_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n316_), .B(new_n318_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n309_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n309_), .B2(new_n324_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT78), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n309_), .A2(new_n324_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n326_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G43gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(G15gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n336_), .B(new_n339_), .Z(new_n340_));
  NAND3_X1  g139(.A1(new_n329_), .A2(new_n334_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n340_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n342_), .B(KEYINPUT78), .C1(new_n327_), .C2(new_n328_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G127gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(G134gat), .ZN(new_n346_));
  INV_X1    g145(.A(G134gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(G127gat), .ZN(new_n348_));
  INV_X1    g147(.A(G113gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(G120gat), .ZN(new_n350_));
  INV_X1    g149(.A(G120gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(G113gat), .ZN(new_n352_));
  OAI22_X1  g151(.A1(new_n346_), .A2(new_n348_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n356_), .A3(KEYINPUT80), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT80), .B1(new_n353_), .B2(new_n356_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT81), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n362_));
  INV_X1    g161(.A(new_n356_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n354_), .A2(new_n355_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n357_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n361_), .A2(new_n368_), .A3(KEYINPUT31), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT79), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT31), .B1(new_n361_), .B2(new_n368_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n344_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n370_), .A2(new_n371_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n280_), .A2(new_n283_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT19), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n290_), .A2(KEYINPUT25), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G183gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n287_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n319_), .A2(new_n321_), .A3(new_n299_), .A4(new_n301_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n323_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n311_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n298_), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n386_), .A2(new_n387_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT20), .B1(new_n391_), .B2(new_n258_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n268_), .B1(new_n309_), .B2(new_n324_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n378_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT89), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n390_), .A2(new_n388_), .ZN(new_n396_));
  AND4_X1   g195(.A1(new_n321_), .A2(new_n319_), .A3(new_n299_), .A4(new_n301_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n385_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n284_), .A2(new_n382_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n287_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n395_), .B1(new_n401_), .B2(new_n268_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n391_), .A2(new_n258_), .A3(KEYINPUT89), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n309_), .A2(new_n268_), .A3(new_n324_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n394_), .B1(new_n405_), .B2(new_n378_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G8gat), .B(G36gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n405_), .A2(new_n378_), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n392_), .A2(new_n393_), .A3(new_n378_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT94), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n412_), .A2(new_n415_), .A3(new_n416_), .A4(KEYINPUT27), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(KEYINPUT27), .A3(new_n415_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT94), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420_));
  INV_X1    g219(.A(new_n415_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n376_), .A2(new_n417_), .A3(new_n419_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n229_), .A2(new_n425_), .A3(new_n365_), .A4(new_n357_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT91), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n360_), .A2(new_n428_), .A3(new_n425_), .A4(new_n229_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT90), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n360_), .A2(new_n229_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n219_), .B(new_n228_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(KEYINPUT4), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G85gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT0), .B(G57gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  INV_X1    g239(.A(new_n432_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n434_), .B(new_n441_), .C1(new_n366_), .C2(new_n231_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT92), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n433_), .A2(new_n444_), .A3(new_n434_), .A4(new_n441_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n436_), .A2(new_n440_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n440_), .B1(new_n436_), .B2(new_n446_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT93), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n436_), .A2(new_n446_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n440_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n447_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n202_), .B1(new_n424_), .B2(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n419_), .A2(new_n417_), .A3(new_n423_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n456_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(KEYINPUT95), .A3(new_n459_), .A4(new_n376_), .ZN(new_n460_));
  AND4_X1   g259(.A1(KEYINPUT33), .A2(new_n436_), .A3(new_n440_), .A4(new_n446_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n433_), .A2(new_n434_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n440_), .B1(new_n462_), .B2(new_n432_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n430_), .A2(new_n441_), .A3(new_n435_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT33), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n461_), .B1(new_n447_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n421_), .A2(new_n422_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n453_), .A2(new_n447_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n410_), .A2(KEYINPUT32), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n404_), .A2(KEYINPUT20), .ZN(new_n471_));
  INV_X1    g270(.A(new_n378_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n403_), .A4(new_n402_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n473_), .B2(new_n394_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n413_), .A2(new_n414_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(new_n470_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n467_), .A2(new_n468_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n280_), .A2(new_n283_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n419_), .A2(new_n417_), .A3(new_n423_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n450_), .A2(new_n455_), .A3(new_n283_), .A4(new_n280_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n477_), .A2(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n373_), .A2(new_n375_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n457_), .A2(new_n460_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G29gat), .B(G36gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G43gat), .B(G50gat), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n486_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G1gat), .A2(G8gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT14), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G1gat), .ZN(new_n496_));
  INV_X1    g295(.A(G8gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n493_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n492_), .A2(new_n493_), .A3(new_n498_), .A4(new_n494_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n487_), .A2(KEYINPUT15), .A3(new_n488_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n491_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n489_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(new_n488_), .A3(new_n487_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n506_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n511_), .A3(KEYINPUT72), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n504_), .A2(new_n513_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G113gat), .B(G141gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(new_n514_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G230gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526_));
  OR2_X1    g325(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n277_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n530_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT65), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT6), .ZN(new_n535_));
  AND2_X1   g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n529_), .B(new_n531_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G85gat), .B(G92gat), .ZN(new_n541_));
  AOI211_X1 g340(.A(new_n530_), .B(new_n540_), .C1(new_n541_), .C2(KEYINPUT9), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n526_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(new_n530_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n541_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n536_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n534_), .A2(KEYINPUT6), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n532_), .A2(KEYINPUT65), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n529_), .A2(new_n531_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n547_), .A2(new_n553_), .A3(new_n554_), .A4(KEYINPUT66), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n543_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557_));
  INV_X1    g356(.A(G99gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n277_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT8), .B1(new_n562_), .B2(new_n541_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n559_), .A2(new_n560_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT8), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n545_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(G78gat), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n265_), .A3(new_n570_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G57gat), .B(G64gat), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n572_), .A2(new_n573_), .B1(KEYINPUT11), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(KEYINPUT11), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n572_), .A2(new_n573_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n575_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n556_), .A2(new_n568_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n556_), .B2(new_n568_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(KEYINPUT68), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n543_), .A2(new_n555_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n578_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n525_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n582_), .B2(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n556_), .A2(new_n568_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n578_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(KEYINPUT12), .A3(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n587_), .A2(new_n590_), .A3(new_n524_), .A4(new_n579_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT5), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n585_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(KEYINPUT13), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n484_), .A2(new_n523_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT34), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n556_), .A2(new_n489_), .A3(new_n568_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n491_), .A2(new_n503_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n556_), .B2(new_n568_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT35), .B(new_n607_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n588_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(KEYINPUT35), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n556_), .A2(new_n568_), .A3(new_n489_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n607_), .A2(KEYINPUT35), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .A4(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT36), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT69), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n621_), .A2(KEYINPUT36), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n611_), .A2(new_n617_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT69), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n618_), .A2(new_n628_), .A3(new_n622_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .A4(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT70), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n625_), .B1(new_n623_), .B2(new_n627_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n630_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n631_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n502_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(new_n578_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT17), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT16), .ZN(new_n643_));
  XOR2_X1   g442(.A(G183gat), .B(G211gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  MUX2_X1   g444(.A(new_n641_), .B(new_n640_), .S(new_n645_), .Z(new_n646_));
  INV_X1    g445(.A(KEYINPUT71), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n639_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n646_), .B(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n636_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n605_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n496_), .A3(new_n456_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT96), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n652_), .A2(new_n655_), .A3(new_n496_), .A4(new_n456_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT97), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n654_), .A2(new_n656_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT38), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(KEYINPUT38), .A3(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n629_), .A2(new_n627_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n628_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT98), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n650_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n605_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G1gat), .B1(new_n671_), .B2(new_n459_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n663_), .A2(new_n664_), .A3(new_n672_), .ZN(G1324gat));
  AOI21_X1  g472(.A(new_n497_), .B1(new_n670_), .B2(new_n479_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT39), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n652_), .A2(new_n497_), .A3(new_n479_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(KEYINPUT40), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1325gat));
  AOI21_X1  g480(.A(new_n338_), .B1(new_n670_), .B2(new_n482_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT41), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n652_), .A2(new_n338_), .A3(new_n482_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n478_), .B(KEYINPUT99), .Z(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n670_), .B2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT42), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n652_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(new_n667_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n649_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n605_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n456_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n604_), .A2(new_n649_), .A3(new_n523_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n665_), .A2(KEYINPUT37), .A3(new_n666_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT70), .B1(new_n697_), .B2(new_n632_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n630_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n484_), .A2(KEYINPUT43), .A3(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT100), .B(KEYINPUT43), .Z(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n457_), .A2(new_n460_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n481_), .A2(new_n483_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n706_), .B2(new_n636_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n696_), .C1(new_n701_), .C2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT101), .ZN(new_n709_));
  INV_X1    g508(.A(new_n696_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n702_), .B1(new_n484_), .B2(new_n700_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n712_), .A3(new_n636_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(KEYINPUT44), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n709_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n696_), .B1(new_n701_), .B2(new_n707_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n456_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n695_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n458_), .A2(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n694_), .B2(new_n725_), .ZN(new_n726_));
  AND4_X1   g525(.A1(new_n724_), .A2(new_n605_), .A3(new_n693_), .A4(new_n725_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n726_), .A2(new_n727_), .B1(KEYINPUT102), .B2(KEYINPUT46), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n717_), .A2(new_n479_), .A3(new_n720_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G36gat), .ZN(new_n730_));
  AND2_X1   g529(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1329gat));
  NAND4_X1  g531(.A1(new_n717_), .A2(G43gat), .A3(new_n482_), .A4(new_n720_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G43gat), .B1(new_n694_), .B2(new_n482_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g536(.A(G50gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n687_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT105), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n694_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n478_), .B1(new_n714_), .B2(KEYINPUT44), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n709_), .B2(new_n716_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n738_), .B1(new_n743_), .B2(KEYINPUT103), .ZN(new_n744_));
  INV_X1    g543(.A(new_n478_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n717_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT104), .B1(new_n744_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n711_), .A2(new_n713_), .ZN(new_n751_));
  AND4_X1   g550(.A1(new_n715_), .A2(new_n751_), .A3(KEYINPUT44), .A4(new_n696_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n715_), .B1(new_n714_), .B2(KEYINPUT44), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n746_), .B(KEYINPUT103), .C1(new_n752_), .C2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G50gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT103), .B1(new_n717_), .B2(new_n746_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n741_), .B1(new_n750_), .B2(new_n758_), .ZN(G1331gat));
  INV_X1    g558(.A(G57gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n706_), .A2(new_n523_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n761_), .A2(KEYINPUT106), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(KEYINPUT106), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n604_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n651_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n760_), .B1(new_n765_), .B2(new_n459_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(KEYINPUT107), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(KEYINPUT107), .ZN(new_n768_));
  AND4_X1   g567(.A1(new_n523_), .A2(new_n706_), .A3(new_n604_), .A4(new_n669_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n459_), .A2(new_n760_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n767_), .A2(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(G1332gat));
  INV_X1    g570(.A(G64gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n769_), .B2(new_n479_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT48), .Z(new_n774_));
  NAND2_X1  g573(.A1(new_n479_), .A2(new_n772_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n765_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT108), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n769_), .B2(new_n482_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT49), .Z(new_n780_));
  NAND2_X1  g579(.A1(new_n482_), .A2(new_n778_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n765_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(G1334gat));
  AOI21_X1  g583(.A(new_n265_), .B1(new_n769_), .B2(new_n687_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT50), .Z(new_n786_));
  NAND2_X1  g585(.A1(new_n687_), .A2(new_n265_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n765_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT110), .ZN(G1335gat));
  NAND4_X1  g588(.A1(new_n762_), .A2(new_n604_), .A3(new_n693_), .A4(new_n763_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(G85gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n456_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n604_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n794_), .A2(new_n522_), .A3(new_n649_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n751_), .A2(new_n795_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n796_), .A2(KEYINPUT111), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(KEYINPUT111), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n459_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n793_), .B1(new_n799_), .B2(new_n792_), .ZN(G1336gat));
  INV_X1    g599(.A(G92gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n790_), .B2(new_n458_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT112), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n798_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n458_), .A2(new_n801_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(G1337gat));
  NAND4_X1  g605(.A1(new_n791_), .A2(new_n527_), .A3(new_n528_), .A4(new_n482_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n483_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n558_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g609(.A(G106gat), .B1(new_n796_), .B2(new_n745_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT52), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n745_), .A2(G106gat), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OR3_X1    g613(.A1(new_n790_), .A2(KEYINPUT113), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT113), .B1(new_n790_), .B2(new_n814_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n812_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n812_), .B2(new_n817_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1339gat));
  AND3_X1   g620(.A1(new_n602_), .A2(new_n523_), .A3(new_n603_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n649_), .C1(new_n635_), .C2(new_n634_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n504_), .A2(new_n510_), .A3(new_n506_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n518_), .B1(new_n509_), .B2(new_n505_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n515_), .A2(new_n518_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n599_), .A2(new_n828_), .ZN(new_n829_));
  AND4_X1   g628(.A1(new_n524_), .A2(new_n587_), .A3(new_n590_), .A4(new_n579_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n579_), .B1(new_n580_), .B2(KEYINPUT12), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n582_), .A2(new_n586_), .A3(new_n578_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n525_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(KEYINPUT55), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n831_), .A2(new_n832_), .A3(new_n835_), .A4(new_n525_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n596_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n829_), .B1(new_n837_), .B2(KEYINPUT56), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n596_), .C1(new_n834_), .C2(new_n836_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT58), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n700_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  INV_X1    g642(.A(new_n829_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n833_), .A2(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n591_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n836_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n598_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n844_), .B1(new_n848_), .B2(new_n839_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n840_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n843_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n636_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n838_), .A2(KEYINPUT58), .A3(new_n840_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n842_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n846_), .A2(new_n847_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n839_), .A4(new_n596_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n837_), .A2(KEYINPUT56), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n837_), .A2(KEYINPUT116), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n599_), .A2(KEYINPUT115), .A3(new_n522_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n599_), .B2(new_n522_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .A4(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n600_), .A2(new_n828_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n692_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT57), .A3(new_n692_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n855_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n825_), .B1(new_n871_), .B2(new_n650_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n424_), .A2(new_n459_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(KEYINPUT118), .Z(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n349_), .A3(new_n522_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(KEYINPUT59), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n523_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n882_), .B2(new_n349_), .ZN(G1340gat));
  OAI21_X1  g682(.A(new_n351_), .B1(new_n794_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n877_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n351_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n794_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n351_), .ZN(G1341gat));
  NAND3_X1  g686(.A1(new_n877_), .A2(new_n345_), .A3(new_n649_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n650_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n345_), .ZN(G1342gat));
  NAND3_X1  g689(.A1(new_n877_), .A2(new_n347_), .A3(new_n668_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n700_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n347_), .ZN(G1343gat));
  NOR4_X1   g692(.A1(new_n459_), .A2(new_n479_), .A3(new_n745_), .A4(new_n482_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n873_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n523_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n214_), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n794_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n215_), .ZN(G1345gat));
  OR3_X1    g698(.A1(new_n895_), .A2(KEYINPUT119), .A3(new_n650_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT119), .B1(new_n895_), .B2(new_n650_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n900_), .A2(new_n901_), .A3(new_n903_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1346gat));
  INV_X1    g706(.A(new_n895_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G162gat), .B1(new_n908_), .B2(new_n668_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n700_), .A2(new_n205_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT120), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n908_), .B2(new_n911_), .ZN(G1347gat));
  INV_X1    g711(.A(new_n687_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n456_), .A2(new_n483_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n479_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n522_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n913_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n918_), .B2(new_n917_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n310_), .B1(new_n873_), .B2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT62), .Z(new_n922_));
  NOR3_X1   g721(.A1(new_n872_), .A2(new_n687_), .A3(new_n915_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(new_n522_), .A3(new_n314_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1348gat));
  AOI21_X1  g724(.A(G176gat), .B1(new_n923_), .B2(new_n604_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n872_), .B2(new_n478_), .ZN(new_n928_));
  AOI21_X1  g727(.A(KEYINPUT57), .B1(new_n866_), .B2(new_n692_), .ZN(new_n929_));
  AOI211_X1 g728(.A(new_n868_), .B(new_n667_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n649_), .B1(new_n931_), .B2(new_n855_), .ZN(new_n932_));
  OAI211_X1 g731(.A(KEYINPUT122), .B(new_n745_), .C1(new_n932_), .C2(new_n825_), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n928_), .A2(new_n916_), .A3(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n794_), .A2(new_n315_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n926_), .B1(new_n934_), .B2(new_n935_), .ZN(G1349gat));
  NAND4_X1  g735(.A1(new_n928_), .A2(new_n649_), .A3(new_n916_), .A4(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n290_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n923_), .B(new_n649_), .C1(new_n385_), .C2(new_n383_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n938_), .A2(KEYINPUT123), .A3(new_n939_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n923_), .A2(new_n287_), .A3(new_n668_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n923_), .A2(new_n636_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n946_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n947_));
  AOI21_X1  g746(.A(KEYINPUT124), .B1(new_n946_), .B2(G190gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n945_), .B1(new_n947_), .B2(new_n948_), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n480_), .A2(new_n482_), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n950_), .B(KEYINPUT125), .Z(new_n951_));
  NOR3_X1   g750(.A1(new_n872_), .A2(new_n458_), .A3(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n522_), .ZN(new_n953_));
  OR3_X1    g752(.A1(new_n953_), .A2(KEYINPUT126), .A3(new_n241_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT126), .B1(new_n953_), .B2(new_n241_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n241_), .ZN(new_n956_));
  AND3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(G1352gat));
  NAND2_X1  g756(.A1(new_n952_), .A2(new_n604_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g758(.A1(new_n952_), .A2(new_n649_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  AND2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n960_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n960_), .B2(new_n961_), .ZN(G1354gat));
  AOI21_X1  g763(.A(G218gat), .B1(new_n952_), .B2(new_n668_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n636_), .A2(G218gat), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(KEYINPUT127), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n965_), .B1(new_n952_), .B2(new_n967_), .ZN(G1355gat));
endmodule


