//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n207_), .B1(KEYINPUT24), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT87), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n207_), .B(KEYINPUT87), .C1(KEYINPUT24), .C2(new_n210_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G169gat), .B(G176gat), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n217_), .B(new_n220_), .C1(new_n221_), .C2(new_n218_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .A4(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT89), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n208_), .A2(new_n209_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT22), .B1(new_n208_), .B2(KEYINPUT88), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n208_), .A2(KEYINPUT22), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n209_), .B(new_n228_), .C1(new_n229_), .C2(KEYINPUT88), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n224_), .A2(KEYINPUT89), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n223_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G197gat), .B(G204gat), .Z(new_n234_));
  INV_X1    g033(.A(KEYINPUT94), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT21), .ZN(new_n236_));
  XOR2_X1   g035(.A(G211gat), .B(G218gat), .Z(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n236_), .A2(new_n237_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n234_), .A2(KEYINPUT21), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n233_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT98), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT22), .B(G169gat), .Z(new_n244_));
  OAI211_X1 g043(.A(new_n224_), .B(new_n227_), .C1(G176gat), .C2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n215_), .A2(new_n246_), .B1(new_n221_), .B2(new_n217_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n247_), .B(new_n207_), .C1(new_n210_), .C2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(new_n241_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT99), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT20), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n243_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT100), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT20), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n249_), .B2(new_n241_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n233_), .B2(new_n241_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n253_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G8gat), .B(G36gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT18), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G64gat), .B(G92gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G155gat), .B(G162gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT92), .ZN(new_n270_));
  INV_X1    g069(.A(G141gat), .ZN(new_n271_));
  INV_X1    g070(.A(G148gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT3), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT2), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(KEYINPUT3), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n270_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G155gat), .ZN(new_n282_));
  INV_X1    g081(.A(G162gat), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT1), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT1), .B1(new_n282_), .B2(new_n283_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n284_), .B(new_n285_), .C1(G155gat), .C2(G162gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(new_n275_), .A3(new_n273_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT93), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G127gat), .B(G134gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT4), .ZN(new_n296_));
  INV_X1    g095(.A(new_n288_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n294_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(KEYINPUT101), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(KEYINPUT101), .B2(new_n295_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n296_), .B1(new_n300_), .B2(KEYINPUT4), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G225gat), .A2(G233gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G29gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G85gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT0), .B(G57gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  INV_X1    g106(.A(new_n302_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n300_), .B2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n266_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n268_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n300_), .A2(new_n308_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n314_), .A2(KEYINPUT33), .A3(new_n307_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT33), .B1(new_n314_), .B2(new_n307_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n314_), .A2(new_n307_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n307_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n266_), .A2(KEYINPUT32), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n257_), .A2(new_n261_), .A3(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n260_), .A2(new_n253_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT102), .ZN(new_n324_));
  INV_X1    g123(.A(new_n243_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n241_), .B(KEYINPUT95), .ZN(new_n326_));
  INV_X1    g125(.A(new_n249_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n258_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n324_), .B1(new_n329_), .B2(new_n254_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT32), .A3(new_n266_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n322_), .A2(new_n331_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n312_), .A2(new_n317_), .B1(new_n320_), .B2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n293_), .B(KEYINPUT31), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT90), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT91), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G15gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n233_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341_));
  INV_X1    g140(.A(G43gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT30), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n340_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT91), .ZN(new_n346_));
  AOI211_X1 g145(.A(new_n337_), .B(new_n345_), .C1(new_n346_), .C2(new_n334_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n345_), .A2(new_n337_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n290_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT28), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G22gat), .B(G50gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n241_), .B(new_n357_), .C1(new_n290_), .C2(new_n351_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n326_), .B1(KEYINPUT29), .B2(new_n288_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n357_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT96), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n360_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n355_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n350_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n366_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n350_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n349_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n318_), .A2(new_n319_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n268_), .B2(new_n311_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n330_), .B2(new_n267_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  OAI22_X1  g177(.A1(new_n333_), .A2(new_n367_), .B1(new_n373_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G230gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G85gat), .ZN(new_n382_));
  INV_X1    g181(.A(G92gat), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n382_), .A2(new_n383_), .A3(KEYINPUT9), .ZN(new_n384_));
  XOR2_X1   g183(.A(G85gat), .B(G92gat), .Z(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(KEYINPUT9), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT10), .B(G99gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT64), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n388_), .B2(G106gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G99gat), .A2(G106gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT6), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(KEYINPUT65), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n390_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n390_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(KEYINPUT65), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(KEYINPUT6), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT66), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(KEYINPUT66), .A3(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n389_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT69), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n395_), .A2(new_n399_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT7), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G99gat), .A2(G106gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(KEYINPUT67), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT67), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n412_), .A2(G99gat), .A3(G106gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT68), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(KEYINPUT67), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n412_), .B1(G99gat), .B2(G106gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .A4(new_n409_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n385_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n406_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n395_), .A2(new_n399_), .A3(new_n407_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(new_n418_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT69), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n425_), .A3(KEYINPUT8), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n402_), .A2(new_n423_), .A3(new_n403_), .A4(new_n407_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT8), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n385_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n405_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G57gat), .B(G64gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G71gat), .B(G78gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n434_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n381_), .B1(new_n430_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT8), .B1(new_n424_), .B2(KEYINPUT69), .ZN(new_n442_));
  AOI211_X1 g241(.A(new_n406_), .B(new_n420_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n429_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n405_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n439_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI211_X1 g247(.A(KEYINPUT12), .B(new_n439_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n440_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n430_), .A2(new_n439_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n444_), .A2(new_n445_), .A3(new_n439_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n381_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G120gat), .B(G148gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT5), .ZN(new_n457_));
  XOR2_X1   g256(.A(G176gat), .B(G204gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT13), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n463_), .B1(KEYINPUT70), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G113gat), .B(G141gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT85), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G169gat), .B(G197gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(G15gat), .B(G22gat), .Z(new_n475_));
  NAND2_X1  g274(.A1(G1gat), .A2(G8gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(KEYINPUT14), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT81), .ZN(new_n478_));
  XOR2_X1   g277(.A(G1gat), .B(G8gat), .Z(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT81), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n477_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n479_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G29gat), .B(G36gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G43gat), .B(G50gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n480_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(KEYINPUT84), .A3(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n474_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n485_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n488_), .B(KEYINPUT15), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n491_), .B(new_n474_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n473_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n473_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n490_), .A2(KEYINPUT84), .A3(new_n491_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT84), .B1(new_n490_), .B2(new_n491_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n500_), .B(new_n503_), .C1(new_n506_), .C2(new_n474_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n469_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n379_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n514_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT35), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n444_), .A2(new_n488_), .A3(new_n445_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n499_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n519_), .B(new_n520_), .C1(new_n521_), .C2(KEYINPUT72), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(KEYINPUT72), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n516_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n515_), .B(KEYINPUT76), .Z(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n430_), .B2(new_n499_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(new_n519_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT77), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n430_), .A2(new_n488_), .B1(new_n518_), .B2(new_n517_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n521_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT77), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .A4(new_n525_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G190gat), .B(G218gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT73), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT74), .B(KEYINPUT75), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n524_), .A2(new_n528_), .A3(new_n532_), .A4(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT78), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n532_), .A2(new_n528_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n524_), .A4(new_n540_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n524_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n536_), .B(KEYINPUT36), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n511_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n551_), .A3(new_n548_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n511_), .A4(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(KEYINPUT79), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n546_), .A2(new_n558_), .A3(new_n511_), .A4(new_n552_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT80), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n550_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT82), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n485_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n439_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT17), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(KEYINPUT17), .A3(new_n570_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n561_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n510_), .A2(new_n575_), .ZN(new_n576_));
  OR3_X1    g375(.A1(new_n576_), .A2(G1gat), .A3(new_n372_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT38), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n555_), .A2(new_n546_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n574_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n510_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(G1gat), .B1(new_n583_), .B2(new_n372_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n578_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n584_), .A3(new_n585_), .ZN(G1324gat));
  INV_X1    g385(.A(new_n378_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G8gat), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n587_), .A2(G8gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n592_));
  OAI221_X1 g391(.A(new_n590_), .B1(new_n576_), .B2(new_n591_), .C1(new_n588_), .C2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(G1325gat));
  OAI21_X1  g394(.A(G15gat), .B1(new_n583_), .B2(new_n350_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT41), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n576_), .A2(G15gat), .A3(new_n350_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(G1326gat));
  XNOR2_X1  g398(.A(new_n368_), .B(KEYINPUT104), .ZN(new_n600_));
  OAI21_X1  g399(.A(G22gat), .B1(new_n583_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT42), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n576_), .A2(G22gat), .A3(new_n600_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT105), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(G1327gat));
  INV_X1    g406(.A(new_n574_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n580_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n510_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(G29gat), .B1(new_n610_), .B2(new_n320_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n509_), .A2(new_n574_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n561_), .B2(KEYINPUT106), .ZN(new_n614_));
  INV_X1    g413(.A(new_n379_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n561_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n379_), .B(new_n561_), .C1(KEYINPUT106), .C2(new_n613_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n612_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT44), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n620_), .A2(G29gat), .A3(new_n320_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(KEYINPUT44), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n611_), .B1(new_n621_), .B2(new_n623_), .ZN(G1328gat));
  INV_X1    g423(.A(G36gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n587_), .B1(new_n619_), .B2(KEYINPUT44), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n587_), .A2(G36gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n610_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(KEYINPUT45), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(KEYINPUT45), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n634_), .A3(KEYINPUT46), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT46), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n627_), .B2(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1329gat));
  NAND2_X1  g437(.A1(new_n610_), .A2(new_n349_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n342_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n620_), .A2(G43gat), .A3(new_n349_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(new_n622_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g442(.A(new_n600_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G50gat), .B1(new_n610_), .B2(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n620_), .A2(G50gat), .A3(new_n368_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n623_), .ZN(G1331gat));
  NAND2_X1  g446(.A1(new_n502_), .A2(new_n507_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n468_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n379_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(new_n575_), .ZN(new_n651_));
  INV_X1    g450(.A(G57gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n320_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n582_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G57gat), .B1(new_n654_), .B2(new_n372_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(G1332gat));
  OAI21_X1  g455(.A(G64gat), .B1(new_n654_), .B2(new_n587_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT107), .Z(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT48), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(KEYINPUT48), .ZN(new_n660_));
  INV_X1    g459(.A(G64gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n651_), .A2(new_n661_), .A3(new_n378_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(G1333gat));
  OAI21_X1  g462(.A(G71gat), .B1(new_n654_), .B2(new_n350_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(G71gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n651_), .A2(new_n667_), .A3(new_n349_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1334gat));
  OAI21_X1  g468(.A(G78gat), .B1(new_n654_), .B2(new_n600_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT50), .ZN(new_n671_));
  INV_X1    g470(.A(G78gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n651_), .A2(new_n672_), .A3(new_n644_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1335gat));
  NAND2_X1  g473(.A1(new_n650_), .A2(new_n609_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n382_), .B1(new_n675_), .B2(new_n372_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT109), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n649_), .A2(new_n574_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT110), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n320_), .A2(G85gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT111), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n677_), .B1(new_n680_), .B2(new_n682_), .ZN(G1336gat));
  AOI21_X1  g482(.A(new_n383_), .B1(new_n680_), .B2(new_n378_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n675_), .A2(G92gat), .A3(new_n587_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1337gat));
  INV_X1    g485(.A(G99gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n680_), .B2(new_n349_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n675_), .A2(new_n388_), .A3(new_n350_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g490(.A(G106gat), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n650_), .A2(new_n692_), .A3(new_n368_), .A4(new_n609_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT52), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n680_), .A2(new_n368_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G106gat), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT52), .B(new_n692_), .C1(new_n680_), .C2(new_n368_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT53), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT53), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n700_), .B(new_n693_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1339gat));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n455_), .A2(new_n459_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n508_), .B2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n460_), .A2(new_n648_), .A3(KEYINPUT113), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n452_), .A2(new_n380_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT12), .B1(new_n430_), .B2(new_n439_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n446_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT114), .B1(new_n711_), .B2(KEYINPUT55), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT114), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT55), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n450_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n440_), .B(KEYINPUT55), .C1(new_n448_), .C2(new_n449_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(KEYINPUT116), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT116), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n711_), .B2(KEYINPUT55), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n712_), .B(new_n715_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n452_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT115), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT115), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n723_), .B(new_n452_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n722_), .A2(new_n724_), .A3(new_n381_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n459_), .B1(new_n720_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n716_), .A2(KEYINPUT116), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n711_), .A2(new_n718_), .A3(KEYINPUT55), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n732_), .A2(new_n725_), .A3(new_n712_), .A4(new_n715_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(KEYINPUT56), .A3(new_n459_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n707_), .B1(new_n729_), .B2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n497_), .A2(new_n499_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n474_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n491_), .A2(new_n737_), .ZN(new_n738_));
  OAI221_X1 g537(.A(new_n473_), .B1(new_n736_), .B2(new_n738_), .C1(new_n506_), .C2(new_n737_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n507_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n463_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT57), .B(new_n580_), .C1(new_n735_), .C2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n557_), .A2(new_n560_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n550_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT58), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT118), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n740_), .A2(new_n704_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n733_), .A2(KEYINPUT56), .A3(new_n459_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT56), .B1(new_n733_), .B2(new_n459_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n746_), .B(new_n747_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n743_), .A2(new_n744_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n729_), .A2(new_n734_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n746_), .B1(new_n752_), .B2(new_n747_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n742_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n580_), .B1(new_n735_), .B2(new_n741_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT117), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n754_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(KEYINPUT117), .A3(new_n756_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n608_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n468_), .A2(new_n508_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n575_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n761_), .ZN(new_n765_));
  NOR4_X1   g564(.A1(new_n561_), .A2(new_n762_), .A3(new_n574_), .A4(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT119), .B1(new_n760_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  INV_X1    g569(.A(new_n706_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT113), .B1(new_n460_), .B2(new_n648_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n741_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n581_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n770_), .B1(new_n776_), .B2(KEYINPUT57), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(KEYINPUT118), .A3(new_n745_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n561_), .A3(new_n750_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n777_), .A2(new_n759_), .A3(new_n742_), .A4(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n574_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n767_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n378_), .A2(new_n372_), .A3(new_n370_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n769_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n648_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n776_), .A2(KEYINPUT57), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n574_), .B1(new_n754_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n767_), .A2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n785_), .A3(new_n793_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n508_), .B(new_n794_), .C1(new_n786_), .C2(KEYINPUT59), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n789_), .B1(new_n795_), .B2(new_n788_), .ZN(G1340gat));
  INV_X1    g595(.A(G120gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n468_), .B2(KEYINPUT60), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n787_), .B(new_n798_), .C1(KEYINPUT60), .C2(new_n797_), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n468_), .B(new_n794_), .C1(new_n786_), .C2(KEYINPUT59), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n797_), .ZN(G1341gat));
  INV_X1    g600(.A(G127gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n787_), .A2(new_n802_), .A3(new_n608_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n574_), .B(new_n794_), .C1(new_n786_), .C2(KEYINPUT59), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n802_), .ZN(G1342gat));
  AOI21_X1  g604(.A(G134gat), .B1(new_n787_), .B2(new_n581_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n794_), .B1(new_n786_), .B2(KEYINPUT59), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT121), .B(G134gat), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n616_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n806_), .B1(new_n807_), .B2(new_n809_), .ZN(G1343gat));
  NAND2_X1  g609(.A1(new_n769_), .A2(new_n784_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n378_), .A2(new_n372_), .A3(new_n369_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n811_), .A2(new_n508_), .A3(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(new_n271_), .ZN(G1344gat));
  NOR3_X1   g614(.A1(new_n811_), .A2(new_n468_), .A3(new_n813_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(new_n272_), .ZN(G1345gat));
  AND3_X1   g616(.A1(new_n782_), .A2(new_n783_), .A3(new_n767_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n783_), .B1(new_n782_), .B2(new_n767_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT61), .B(G155gat), .Z(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n820_), .A2(new_n608_), .A3(new_n812_), .A4(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n769_), .A2(new_n608_), .A3(new_n784_), .A4(new_n812_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n821_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n823_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1346gat));
  NAND4_X1  g628(.A1(new_n820_), .A2(new_n283_), .A3(new_n581_), .A4(new_n812_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n811_), .A2(new_n616_), .A3(new_n813_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n283_), .ZN(G1347gat));
  NOR2_X1   g631(.A1(new_n587_), .A2(new_n320_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n349_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n644_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n792_), .A2(new_n835_), .ZN(new_n836_));
  OR3_X1    g635(.A1(new_n836_), .A2(KEYINPUT124), .A3(new_n508_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT124), .B1(new_n836_), .B2(new_n508_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(G169gat), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n837_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n838_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n836_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n648_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n841_), .B(new_n842_), .C1(new_n244_), .C2(new_n844_), .ZN(G1348gat));
  AOI21_X1  g644(.A(G176gat), .B1(new_n843_), .B2(new_n469_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n811_), .A2(new_n368_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n834_), .A2(new_n209_), .A3(new_n468_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(G1349gat));
  NOR3_X1   g648(.A1(new_n836_), .A2(new_n217_), .A3(new_n574_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n847_), .A2(new_n349_), .A3(new_n608_), .A4(new_n833_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n203_), .ZN(G1350gat));
  OAI21_X1  g651(.A(G190gat), .B1(new_n836_), .B2(new_n616_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n581_), .A2(new_n221_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT125), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n836_), .B2(new_n855_), .ZN(G1351gat));
  INV_X1    g655(.A(new_n833_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n369_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n820_), .A2(new_n648_), .A3(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT126), .B(G197gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1352gat));
  INV_X1    g660(.A(new_n858_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n811_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n469_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT127), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(G204gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT127), .B(G204gat), .Z(new_n867_));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n469_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1353gat));
  NAND3_X1  g668(.A1(new_n820_), .A2(new_n608_), .A3(new_n858_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT63), .B(G211gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n870_), .B2(new_n873_), .ZN(G1354gat));
  INV_X1    g673(.A(G218gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n863_), .A2(new_n875_), .A3(new_n581_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n811_), .A2(new_n616_), .A3(new_n862_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(new_n877_), .ZN(G1355gat));
endmodule


