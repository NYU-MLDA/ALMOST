//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_;
  NOR2_X1   g000(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n206_));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(KEYINPUT64), .B2(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n221_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n213_), .A2(new_n222_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT66), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n232_), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n233_), .B2(KEYINPUT66), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT66), .B1(new_n229_), .B2(KEYINPUT67), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT7), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n213_), .A2(new_n230_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n216_), .A2(new_n219_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n228_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT65), .B(KEYINPUT6), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n212_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n230_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(new_n236_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n228_), .B(new_n238_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n210_), .B(new_n227_), .C1(new_n239_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT12), .ZN(new_n248_));
  INV_X1    g047(.A(new_n227_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n238_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT8), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n251_), .B2(new_n245_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(new_n210_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n227_), .B1(new_n239_), .B2(new_n246_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  INV_X1    g055(.A(new_n210_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n203_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n257_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n247_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n203_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n252_), .A2(KEYINPUT68), .A3(new_n210_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT5), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G176gat), .B(G204gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  NOR2_X1   g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n267_), .A2(new_n271_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n202_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n279_), .B(KEYINPUT70), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT37), .ZN(new_n282_));
  XOR2_X1   g081(.A(G190gat), .B(G218gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(G134gat), .B(G162gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G29gat), .B(G36gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G43gat), .B(G50gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n291_), .A2(new_n292_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT35), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G232gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT34), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n252_), .A2(new_n296_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n289_), .B(KEYINPUT71), .ZN(new_n302_));
  INV_X1    g101(.A(new_n292_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(new_n293_), .A3(KEYINPUT15), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT15), .B1(new_n304_), .B2(new_n293_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n308_), .A2(new_n252_), .A3(KEYINPUT72), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n310_));
  INV_X1    g109(.A(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n305_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n255_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n301_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n300_), .A2(new_n297_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n317_), .B(new_n301_), .C1(new_n309_), .C2(new_n313_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n288_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n282_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n318_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT72), .B1(new_n308_), .B2(new_n252_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n255_), .A2(new_n312_), .A3(new_n310_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n317_), .B1(new_n325_), .B2(new_n301_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n287_), .B1(new_n322_), .B2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n285_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT74), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n316_), .A2(new_n318_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(KEYINPUT76), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n321_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n321_), .B2(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n331_), .ZN(new_n337_));
  OAI22_X1  g136(.A1(new_n335_), .A2(new_n336_), .B1(KEYINPUT37), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G15gat), .B(G22gat), .ZN(new_n339_));
  INV_X1    g138(.A(G1gat), .ZN(new_n340_));
  INV_X1    g139(.A(G8gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT14), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G8gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(new_n210_), .Z(new_n346_));
  NAND2_X1  g145(.A1(G231gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G127gat), .B(G155gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(G183gat), .B(G211gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n349_), .A2(KEYINPUT17), .A3(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(KEYINPUT17), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n338_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n281_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362_));
  INV_X1    g161(.A(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(G15gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n364_), .B(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT24), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G190gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT26), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT26), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G190gat), .ZN(new_n379_));
  INV_X1    g178(.A(G183gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT25), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G183gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n377_), .A2(new_n379_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n372_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT24), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n384_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n388_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n375_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n376_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n371_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n394_));
  OR3_X1    g193(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n368_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n399_), .A2(new_n400_), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  XNOR2_X1  g202(.A(G113gat), .B(G120gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G134gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G127gat), .ZN(new_n407_));
  INV_X1    g206(.A(G127gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G134gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(KEYINPUT83), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT83), .B1(new_n407_), .B2(new_n409_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n405_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n409_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n410_), .A3(new_n404_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT31), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n403_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n403_), .A2(new_n419_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G197gat), .B(G204gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT21), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G218gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G211gat), .ZN(new_n435_));
  INV_X1    g234(.A(G211gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G218gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G197gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G204gat), .ZN(new_n440_));
  INV_X1    g239(.A(G204gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G197gat), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT86), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT21), .B1(new_n440_), .B2(KEYINPUT86), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n433_), .B(new_n438_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n432_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n435_), .A2(new_n437_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n446_), .A2(KEYINPUT87), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT87), .B1(new_n446_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n445_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT88), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n445_), .B(new_n452_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n396_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n384_), .A2(new_n387_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT80), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n384_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n455_), .B1(new_n459_), .B2(new_n375_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n430_), .B1(new_n454_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n386_), .B(KEYINPUT94), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT22), .B(G169gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT95), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n393_), .B(new_n462_), .C1(new_n465_), .C2(G176gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n381_), .A2(new_n383_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n377_), .A2(new_n379_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n381_), .A2(new_n383_), .A3(KEYINPUT90), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT91), .B1(new_n386_), .B2(KEYINPUT24), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n372_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n386_), .A2(KEYINPUT91), .A3(KEYINPUT24), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(new_n476_), .A3(KEYINPUT92), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n371_), .A2(KEYINPUT93), .A3(new_n374_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT93), .B1(new_n371_), .B2(new_n374_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT92), .B1(new_n472_), .B2(new_n476_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n466_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n450_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n429_), .B1(new_n461_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n397_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n443_), .A2(new_n444_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n447_), .B1(new_n432_), .B2(new_n431_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n441_), .A2(G197gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n439_), .A2(G204gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT21), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n492_), .B2(new_n438_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n446_), .A2(KEYINPUT87), .A3(new_n447_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n487_), .A2(new_n488_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n495_), .B(new_n466_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n486_), .A2(new_n496_), .A3(KEYINPUT20), .A4(new_n429_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G8gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n485_), .A2(new_n498_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n453_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n493_), .A2(new_n494_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n452_), .B1(new_n507_), .B2(new_n445_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n460_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT20), .ZN(new_n510_));
  INV_X1    g309(.A(new_n482_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n495_), .B1(new_n512_), .B2(new_n466_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n428_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n505_), .B1(new_n514_), .B2(new_n497_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n425_), .B1(new_n504_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT29), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G155gat), .A2(G162gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT1), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT1), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(G155gat), .A3(G162gat), .ZN(new_n521_));
  OR2_X1    g320(.A1(G155gat), .A2(G162gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G141gat), .A2(G148gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G141gat), .A2(G148gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT84), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT84), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT3), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT2), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT85), .B1(new_n526_), .B2(new_n533_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT85), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n540_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n522_), .A2(new_n518_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n517_), .B1(new_n532_), .B2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(G228gat), .B(G233gat), .C1(new_n547_), .C2(new_n495_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n523_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n530_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n544_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT29), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G228gat), .A2(G233gat), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n451_), .A3(new_n554_), .A4(new_n453_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G78gat), .B(G106gat), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n532_), .A2(new_n546_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT28), .B1(new_n559_), .B2(KEYINPUT29), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n552_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n517_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G22gat), .B(G50gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n559_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n562_), .B1(new_n561_), .B2(new_n517_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n564_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n557_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n548_), .A2(new_n555_), .A3(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n558_), .A2(new_n566_), .A3(new_n569_), .A4(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n566_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n548_), .A2(new_n570_), .A3(new_n555_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n570_), .B1(new_n548_), .B2(new_n555_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G29gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(G85gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT0), .B(G57gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  OAI21_X1  g380(.A(new_n418_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n532_), .A2(new_n546_), .A3(new_n417_), .A4(new_n413_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G225gat), .A2(G233gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n581_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT4), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT4), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n589_), .B(new_n418_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n586_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT97), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n590_), .A2(new_n586_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT4), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n587_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n588_), .A2(KEYINPUT97), .A3(new_n591_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n599_));
  OAI22_X1  g398(.A1(new_n598_), .A2(new_n599_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n581_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n486_), .A2(new_n496_), .A3(KEYINPUT20), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n428_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n484_), .A2(KEYINPUT20), .A3(new_n509_), .A4(new_n429_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n503_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n514_), .A2(new_n497_), .A3(new_n505_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(KEYINPUT27), .A3(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n516_), .A2(new_n577_), .A3(new_n602_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n572_), .A2(new_n576_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n587_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n614_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n584_), .A2(new_n586_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n617_), .B2(new_n581_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(KEYINPUT102), .A3(new_n516_), .A4(new_n609_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n612_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n590_), .A2(new_n585_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n588_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n582_), .A2(new_n583_), .A3(new_n586_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n601_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n595_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n628_), .A2(KEYINPUT99), .A3(new_n601_), .A4(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n503_), .B1(new_n485_), .B2(new_n498_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(new_n608_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n597_), .A2(KEYINPUT33), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT98), .B1(new_n597_), .B2(KEYINPUT33), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n615_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .A4(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n505_), .A2(KEYINPUT32), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n514_), .A2(new_n497_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n514_), .A2(KEYINPUT100), .A3(new_n497_), .A4(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n639_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n618_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n577_), .B1(new_n638_), .B2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT103), .B(new_n423_), .C1(new_n621_), .C2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n516_), .A2(new_n609_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n422_), .A2(new_n613_), .A3(new_n602_), .A4(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n634_), .A2(new_n637_), .ZN(new_n653_));
  AND4_X1   g452(.A1(new_n633_), .A2(new_n630_), .A3(new_n608_), .A4(new_n631_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n602_), .A2(new_n645_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n653_), .A2(new_n654_), .B1(new_n655_), .B2(new_n644_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n612_), .B(new_n620_), .C1(new_n656_), .C2(new_n577_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT103), .B1(new_n657_), .B2(new_n423_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n652_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT79), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n345_), .A2(new_n293_), .A3(new_n304_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(G229gat), .A2(G233gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n345_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n312_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n662_), .B1(new_n666_), .B2(new_n661_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G113gat), .B(G141gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(G169gat), .B(G197gat), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n669_), .B(new_n670_), .Z(new_n671_));
  AOI21_X1  g470(.A(new_n660_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  NOR4_X1   g472(.A1(new_n665_), .A2(new_n667_), .A3(KEYINPUT79), .A4(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n668_), .A2(new_n671_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n659_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n361_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n602_), .A2(KEYINPUT104), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n602_), .A2(KEYINPUT104), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n340_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT38), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n659_), .A2(new_n337_), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n677_), .B(new_n358_), .C1(new_n276_), .C2(new_n278_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G1gat), .B1(new_n691_), .B2(new_n602_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n686_), .A2(new_n687_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(new_n692_), .A3(new_n693_), .ZN(G1324gat));
  INV_X1    g493(.A(new_n650_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n341_), .A3(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n689_), .A2(new_n695_), .A3(new_n690_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT39), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(G8gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n697_), .B2(G8gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n702_), .B(new_n704_), .ZN(G1325gat));
  OAI21_X1  g504(.A(G15gat), .B1(new_n691_), .B2(new_n423_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT41), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n681_), .A2(new_n366_), .A3(new_n422_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1326gat));
  OAI21_X1  g508(.A(G22gat), .B1(new_n691_), .B2(new_n613_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT42), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n613_), .A2(G22gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n680_), .B2(new_n712_), .ZN(G1327gat));
  NOR2_X1   g512(.A1(new_n337_), .A2(new_n359_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n279_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n659_), .A2(new_n678_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT109), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n659_), .A2(new_n718_), .A3(new_n678_), .A4(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  OR3_X1    g519(.A1(new_n720_), .A2(G29gat), .A3(new_n602_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n279_), .A2(new_n678_), .A3(new_n358_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT106), .Z(new_n723_));
  NOR2_X1   g522(.A1(new_n337_), .A2(KEYINPUT37), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n321_), .A2(new_n332_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT77), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n726_), .B2(new_n334_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n652_), .B2(new_n658_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(KEYINPUT43), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n728_), .B2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n723_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(KEYINPUT44), .B(new_n723_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n685_), .A3(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT108), .B1(new_n736_), .B2(G29gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n721_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  NAND3_X1  g538(.A1(new_n734_), .A2(new_n695_), .A3(new_n735_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G36gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n650_), .A2(G36gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n717_), .A2(new_n719_), .A3(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n741_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(KEYINPUT46), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n741_), .B(new_n745_), .C1(new_n747_), .C2(KEYINPUT46), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1329gat));
  NAND4_X1  g550(.A1(new_n734_), .A2(G43gat), .A3(new_n422_), .A4(new_n735_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n363_), .B1(new_n720_), .B2(new_n423_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g554(.A1(new_n734_), .A2(G50gat), .A3(new_n577_), .A4(new_n735_), .ZN(new_n756_));
  INV_X1    g555(.A(G50gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n720_), .B2(new_n613_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1331gat));
  NAND2_X1  g558(.A1(new_n359_), .A2(new_n677_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n280_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n689_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n602_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n659_), .A2(new_n677_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n360_), .A2(new_n279_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n684_), .A2(G57gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1332gat));
  INV_X1    g567(.A(new_n766_), .ZN(new_n769_));
  INV_X1    g568(.A(G64gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n695_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n762_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n772_), .B2(new_n695_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n773_), .A2(new_n774_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n771_), .B1(new_n776_), .B2(new_n777_), .ZN(G1333gat));
  INV_X1    g577(.A(G71gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n769_), .A2(new_n779_), .A3(new_n422_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n772_), .B2(new_n422_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n781_), .A2(new_n782_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n784_), .B2(new_n785_), .ZN(G1334gat));
  INV_X1    g585(.A(G78gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n769_), .A2(new_n787_), .A3(new_n577_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n772_), .B2(new_n577_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n789_), .A2(new_n790_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n788_), .B1(new_n792_), .B2(new_n793_), .ZN(G1335gat));
  NAND3_X1  g593(.A1(new_n764_), .A2(new_n281_), .A3(new_n714_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n214_), .A3(new_n685_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n730_), .A2(new_n731_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n279_), .A2(new_n678_), .A3(new_n359_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n618_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n797_), .B1(new_n802_), .B2(new_n214_), .ZN(G1336gat));
  OAI21_X1  g602(.A(new_n215_), .B1(new_n795_), .B2(new_n650_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT112), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n650_), .A2(new_n215_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n800_), .B2(new_n806_), .ZN(G1337gat));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n422_), .B(new_n799_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(G99gat), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n422_), .A2(new_n223_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812_));
  OAI22_X1  g611(.A1(new_n795_), .A2(new_n811_), .B1(KEYINPUT114), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(KEYINPUT114), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n809_), .A2(new_n808_), .A3(G99gat), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1338gat));
  NAND3_X1  g618(.A1(new_n796_), .A2(new_n224_), .A3(new_n577_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n577_), .B(new_n799_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(G106gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n821_), .B2(G106gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g625(.A(new_n760_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n338_), .B(new_n827_), .C1(KEYINPUT115), .C2(KEYINPUT54), .ZN(new_n828_));
  NOR2_X1   g627(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n829_));
  INV_X1    g628(.A(new_n278_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n677_), .B(new_n359_), .C1(new_n830_), .C2(new_n275_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n727_), .B2(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n828_), .A2(new_n832_), .B1(KEYINPUT115), .B2(KEYINPUT54), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n666_), .A2(new_n661_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n662_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n308_), .A2(new_n345_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n661_), .A2(new_n835_), .ZN(new_n837_));
  OAI221_X1 g636(.A(new_n673_), .B1(new_n834_), .B2(new_n835_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT118), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n841_), .B(new_n838_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n274_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n272_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n677_), .A2(new_n272_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n260_), .A2(KEYINPUT116), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n256_), .B1(new_n252_), .B2(new_n210_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n261_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n264_), .B1(new_n851_), .B2(new_n258_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(new_n852_), .B2(KEYINPUT55), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT55), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n264_), .A3(new_n258_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n848_), .A2(new_n853_), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT117), .B1(new_n856_), .B2(new_n271_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n846_), .B1(new_n857_), .B2(KEYINPUT56), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n859_));
  AOI211_X1 g658(.A(KEYINPUT117), .B(new_n859_), .C1(new_n856_), .C2(new_n271_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n845_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n337_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(KEYINPUT57), .A3(new_n337_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n272_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n856_), .A2(new_n859_), .A3(new_n271_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n859_), .B1(new_n856_), .B2(new_n271_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n870_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n872_), .A2(KEYINPUT58), .A3(new_n868_), .A4(new_n867_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n727_), .A2(new_n871_), .A3(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n864_), .A2(new_n865_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n833_), .B1(new_n875_), .B2(new_n358_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n422_), .A2(new_n613_), .A3(new_n650_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n684_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(G113gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n881_), .A3(new_n678_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n878_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n876_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n883_), .B2(KEYINPUT119), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n861_), .B2(new_n337_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n727_), .A2(new_n871_), .A3(new_n873_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n359_), .B1(new_n891_), .B2(new_n865_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n878_), .B(new_n888_), .C1(new_n892_), .C2(new_n833_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n887_), .A2(KEYINPUT121), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(KEYINPUT121), .B1(new_n887_), .B2(new_n893_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n677_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n882_), .B1(new_n896_), .B2(new_n881_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n279_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n880_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n280_), .B1(new_n887_), .B2(new_n893_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n898_), .ZN(G1341gat));
  NAND3_X1  g701(.A1(new_n880_), .A2(new_n408_), .A3(new_n359_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n894_), .A2(new_n895_), .A3(new_n358_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n408_), .ZN(G1342gat));
  NOR3_X1   g704(.A1(new_n876_), .A2(new_n337_), .A3(new_n879_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(KEYINPUT122), .A3(new_n406_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n906_), .B2(G134gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n894_), .A2(new_n895_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n338_), .A2(new_n406_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1343gat));
  INV_X1    g713(.A(new_n876_), .ZN(new_n915_));
  NOR4_X1   g714(.A1(new_n422_), .A2(new_n695_), .A3(new_n684_), .A4(new_n613_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n678_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n281_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g721(.A1(new_n917_), .A2(new_n358_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT61), .B(G155gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1346gat));
  OR3_X1    g724(.A1(new_n917_), .A2(G162gat), .A3(new_n337_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G162gat), .B1(new_n917_), .B2(new_n338_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1347gat));
  NOR3_X1   g727(.A1(new_n423_), .A2(new_n650_), .A3(new_n685_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n678_), .ZN(new_n930_));
  OR3_X1    g729(.A1(new_n876_), .A2(new_n577_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(new_n932_), .A3(G169gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n876_), .A2(new_n577_), .A3(new_n930_), .ZN(new_n934_));
  INV_X1    g733(.A(G169gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(KEYINPUT123), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n933_), .A2(KEYINPUT62), .A3(new_n936_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n931_), .A2(new_n465_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n937_), .B(new_n938_), .C1(KEYINPUT62), .C2(new_n936_), .ZN(G1348gat));
  NAND3_X1  g738(.A1(new_n915_), .A2(new_n613_), .A3(new_n929_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G176gat), .B1(new_n940_), .B2(new_n280_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n279_), .A2(G176gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1349gat));
  AND2_X1   g742(.A1(new_n469_), .A2(new_n471_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n940_), .A2(new_n358_), .ZN(new_n945_));
  MUX2_X1   g744(.A(G183gat), .B(new_n944_), .S(new_n945_), .Z(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n940_), .B2(new_n338_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n327_), .A2(new_n470_), .A3(new_n331_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n940_), .B2(new_n948_), .ZN(G1351gat));
  NOR4_X1   g748(.A1(new_n422_), .A2(new_n613_), .A3(new_n618_), .A4(new_n650_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n915_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n677_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(new_n439_), .ZN(G1352gat));
  NOR2_X1   g752(.A1(new_n951_), .A2(new_n280_), .ZN(new_n954_));
  XOR2_X1   g753(.A(KEYINPUT124), .B(G204gat), .Z(new_n955_));
  XNOR2_X1  g754(.A(new_n954_), .B(new_n955_), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n915_), .A2(new_n359_), .A3(new_n950_), .ZN(new_n957_));
  XOR2_X1   g756(.A(KEYINPUT63), .B(G211gat), .Z(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  OAI21_X1  g758(.A(KEYINPUT125), .B1(new_n957_), .B2(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT63), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n957_), .A2(new_n961_), .A3(new_n436_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n962_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n957_), .A2(KEYINPUT125), .A3(new_n959_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1354gat));
  NOR2_X1   g764(.A1(new_n338_), .A2(new_n434_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(KEYINPUT127), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n951_), .A2(new_n967_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n951_), .A2(KEYINPUT126), .A3(new_n337_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(G218gat), .ZN(new_n970_));
  OAI21_X1  g769(.A(KEYINPUT126), .B1(new_n951_), .B2(new_n337_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n968_), .B1(new_n970_), .B2(new_n971_), .ZN(G1355gat));
endmodule


