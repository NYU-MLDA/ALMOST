//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT79), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G71gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G99gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT75), .B(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207_));
  OR3_X1    g006(.A1(new_n206_), .A2(KEYINPUT76), .A3(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(G183gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT76), .B1(new_n206_), .B2(new_n207_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n217_), .B(new_n218_), .C1(new_n221_), .C2(KEYINPUT24), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT77), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G169gat), .A3(G176gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(KEYINPUT24), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n222_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n226_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n206_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n216_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n217_), .A2(new_n218_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n231_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n219_), .A2(KEYINPUT22), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  AOI21_X1  g036(.A(G176gat), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT22), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G169gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n241_), .B2(new_n237_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n213_), .A2(new_n230_), .B1(new_n235_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n205_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT81), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n244_), .A2(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT80), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT30), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT31), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n250_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT82), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(G155gat), .A3(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n260_), .B1(new_n265_), .B2(KEYINPUT1), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(new_n264_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT83), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n262_), .A2(new_n264_), .A3(KEYINPUT83), .A4(new_n267_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G141gat), .B(G148gat), .Z(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n278_), .A2(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(KEYINPUT84), .B2(new_n278_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  OR3_X1    g080(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n260_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n274_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n248_), .A2(new_n286_), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n287_), .A2(KEYINPUT96), .A3(KEYINPUT4), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n272_), .A2(new_n273_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n249_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(KEYINPUT4), .A3(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT96), .B1(new_n287_), .B2(KEYINPUT4), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n288_), .A2(new_n291_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G1gat), .B(G29gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(G57gat), .B(G85gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n290_), .A2(new_n287_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n292_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n295_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(KEYINPUT33), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n295_), .A2(KEYINPUT33), .A3(new_n300_), .A4(new_n302_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n301_), .B2(new_n293_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n288_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n293_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT19), .ZN(new_n310_));
  INV_X1    g109(.A(G218gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G211gat), .ZN(new_n312_));
  INV_X1    g111(.A(G211gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G218gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n316_));
  INV_X1    g115(.A(G197gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G204gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n322_), .B1(G197gat), .B2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n315_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT88), .B1(new_n317_), .B2(G204gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT88), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n319_), .A3(G197gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n318_), .A2(G204gat), .A3(new_n320_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n322_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT89), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n322_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n333_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n331_), .B(new_n332_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n328_), .A2(new_n329_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT89), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n332_), .B1(new_n342_), .B2(new_n331_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n243_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT20), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n331_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n236_), .A2(new_n240_), .A3(new_n220_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT94), .B1(new_n348_), .B2(new_n231_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT94), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n236_), .A2(new_n240_), .A3(new_n220_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n227_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n215_), .A2(new_n216_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n217_), .A2(new_n218_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT95), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n353_), .A2(new_n359_), .A3(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n215_), .A2(KEYINPUT25), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n211_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(new_n221_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n223_), .A3(new_n221_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n363_), .A2(new_n234_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n347_), .B1(new_n361_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n310_), .B1(new_n345_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT18), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  NAND2_X1  g172(.A1(new_n346_), .A2(KEYINPUT90), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n213_), .A2(new_n230_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n235_), .A2(new_n242_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n374_), .B(new_n338_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n359_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n378_));
  AOI211_X1 g177(.A(KEYINPUT95), .B(new_n355_), .C1(new_n349_), .C2(new_n352_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n347_), .B(new_n367_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n310_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n369_), .A2(new_n373_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n373_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n310_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n374_), .A2(new_n338_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n381_), .B1(new_n387_), .B2(new_n243_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n367_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n346_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n383_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n385_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n305_), .A2(new_n308_), .A3(new_n384_), .A4(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n300_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n303_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n387_), .A2(new_n243_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n357_), .A2(new_n367_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT20), .B1(new_n399_), .B2(new_n346_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n310_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n391_), .A2(new_n392_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n404_));
  MUX2_X1   g203(.A(new_n402_), .B(new_n403_), .S(new_n404_), .Z(new_n405_));
  OAI22_X1  g204(.A1(new_n304_), .A2(new_n394_), .B1(new_n396_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n407_), .A2(new_n374_), .A3(new_n338_), .A4(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n346_), .B1(new_n289_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n408_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT91), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(G50gat), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n286_), .A2(KEYINPUT29), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n289_), .B2(new_n412_), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT28), .B(G22gat), .Z(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n419_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n418_), .B1(new_n286_), .B2(KEYINPUT29), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n289_), .A2(new_n412_), .A3(new_n420_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n422_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n417_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n417_), .B2(new_n428_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n409_), .A2(new_n415_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n410_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n416_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n430_), .A2(new_n431_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n434_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n374_), .A2(new_n338_), .A3(new_n408_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n438_), .A2(new_n407_), .B1(new_n414_), .B2(new_n413_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n439_), .B2(new_n411_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n427_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n425_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT92), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n417_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n436_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n435_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n406_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n434_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n436_), .A3(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT27), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n373_), .B1(new_n369_), .B2(new_n383_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n391_), .A2(new_n392_), .A3(new_n385_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n402_), .A2(new_n385_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT27), .A3(new_n384_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n451_), .A2(new_n396_), .A3(new_n455_), .A4(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n259_), .B1(new_n448_), .B2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n373_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n454_), .A2(new_n460_), .A3(new_n452_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT27), .B1(new_n384_), .B2(new_n393_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT98), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT98), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n447_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT98), .B1(new_n461_), .B2(new_n462_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n455_), .A2(new_n464_), .A3(new_n457_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT99), .A3(new_n447_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n259_), .A2(new_n396_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n459_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT71), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G43gat), .B(G50gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G8gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n477_), .A2(KEYINPUT71), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n477_), .A2(KEYINPUT71), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n479_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n481_), .A2(new_n488_), .A3(new_n489_), .A4(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496_));
  INV_X1    g295(.A(new_n492_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n479_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n481_), .A2(KEYINPUT15), .A3(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(new_n488_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n495_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n481_), .A2(new_n492_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n502_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n494_), .B1(new_n505_), .B2(new_n493_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n503_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n497_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT15), .B1(new_n481_), .B2(new_n492_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n502_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n495_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n506_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n509_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n511_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT10), .B(G99gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT64), .B(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(KEYINPUT9), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n524_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G85gat), .ZN(new_n530_));
  INV_X1    g329(.A(G92gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(KEYINPUT9), .A3(new_n523_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT66), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n526_), .A2(new_n528_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n537_));
  OR3_X1    g336(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n523_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT8), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n540_), .B2(KEYINPUT65), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(new_n544_), .A3(new_n541_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n522_), .A2(new_n529_), .A3(new_n548_), .A4(new_n533_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n535_), .A2(new_n546_), .A3(new_n547_), .A4(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n501_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n546_), .A2(new_n547_), .A3(new_n534_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(new_n504_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT35), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(KEYINPUT73), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT72), .ZN(new_n561_));
  XOR2_X1   g360(.A(G134gat), .B(G162gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n551_), .A2(new_n553_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n556_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n558_), .B(KEYINPUT73), .C1(new_n567_), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT74), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n570_), .B(new_n566_), .C1(KEYINPUT36), .C2(new_n564_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n581_));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n502_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(KEYINPUT17), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .A4(KEYINPUT37), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n578_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n546_), .A2(new_n547_), .A3(new_n534_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n585_), .ZN(new_n605_));
  INV_X1    g404(.A(G230gat), .ZN(new_n606_));
  INV_X1    g405(.A(G233gat), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n585_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n583_), .A2(KEYINPUT12), .A3(new_n584_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n550_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n605_), .A2(new_n609_), .A3(new_n610_), .A4(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n604_), .A2(new_n585_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n585_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n552_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n608_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT68), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n602_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n614_), .A2(new_n625_), .A3(new_n618_), .A4(KEYINPUT69), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n619_), .A2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT13), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(KEYINPUT13), .A3(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n601_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n476_), .A2(new_n519_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n396_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n483_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n573_), .A2(new_n575_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n476_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n519_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n633_), .A2(new_n646_), .A3(new_n634_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n633_), .A2(KEYINPUT100), .A3(new_n646_), .A4(new_n634_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n645_), .A2(new_n599_), .A3(new_n649_), .A4(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n396_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n640_), .A2(new_n641_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n642_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT101), .Z(G1324gat));
  XNOR2_X1  g454(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658_));
  INV_X1    g457(.A(new_n471_), .ZN(new_n659_));
  AND4_X1   g458(.A1(new_n659_), .A2(new_n649_), .A3(new_n599_), .A4(new_n650_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n474_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n643_), .B(new_n660_), .C1(new_n661_), .C2(new_n459_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n662_), .A2(new_n663_), .A3(G8gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n662_), .B2(G8gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT39), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(G8gat), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT102), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n662_), .A2(new_n663_), .A3(G8gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n638_), .A2(new_n484_), .A3(new_n659_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n658_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT104), .B(new_n673_), .C1(new_n666_), .C2(new_n671_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n657_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n664_), .A2(new_n665_), .A3(KEYINPUT39), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n669_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n674_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT104), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n672_), .A2(new_n658_), .A3(new_n674_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n656_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n677_), .A2(new_n683_), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n638_), .A2(new_n685_), .A3(new_n259_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT105), .Z(new_n687_));
  INV_X1    g486(.A(new_n259_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G15gat), .B1(new_n651_), .B2(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n689_), .A2(KEYINPUT41), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(KEYINPUT41), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n687_), .A2(new_n690_), .A3(new_n691_), .ZN(G1326gat));
  OAI21_X1  g491(.A(G22gat), .B1(new_n651_), .B2(new_n447_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT42), .ZN(new_n694_));
  INV_X1    g493(.A(G22gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n638_), .A2(new_n695_), .A3(new_n451_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n476_), .A2(new_n519_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n644_), .A2(new_n598_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n635_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n701_), .A2(G29gat), .A3(new_n396_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n578_), .A2(new_n600_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n476_), .B2(new_n704_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n471_), .A2(KEYINPUT99), .A3(new_n447_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT99), .B1(new_n471_), .B2(new_n447_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n475_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n459_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n703_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n705_), .A2(new_n712_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n649_), .A2(new_n598_), .A3(new_n650_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n714_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(KEYINPUT106), .A3(new_n639_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G29gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT106), .B1(new_n718_), .B2(new_n639_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n702_), .B1(new_n720_), .B2(new_n721_), .ZN(G1328gat));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n713_), .A2(new_n714_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n659_), .A3(new_n715_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n701_), .A2(G36gat), .A3(new_n471_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT45), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n723_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n730_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n727_), .A2(G36gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1329gat));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(G43gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n718_), .B2(new_n259_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n259_), .A2(new_n737_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n701_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n716_), .A2(new_n717_), .A3(new_n688_), .ZN(new_n742_));
  OAI221_X1 g541(.A(KEYINPUT47), .B1(new_n701_), .B2(new_n739_), .C1(new_n742_), .C2(new_n737_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1330gat));
  INV_X1    g543(.A(new_n701_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G50gat), .B1(new_n745_), .B2(new_n451_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n451_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n718_), .B2(new_n747_), .ZN(G1331gat));
  NAND4_X1  g547(.A1(new_n645_), .A2(new_n519_), .A3(new_n635_), .A4(new_n599_), .ZN(new_n749_));
  INV_X1    g548(.A(G57gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT110), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n750_), .A2(KEYINPUT110), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n396_), .B(new_n749_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n635_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n601_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT107), .Z(new_n756_));
  NOR2_X1   g555(.A1(new_n476_), .A2(new_n646_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT108), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n750_), .B1(new_n759_), .B2(new_n396_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n760_), .A2(KEYINPUT109), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(KEYINPUT109), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n753_), .B1(new_n761_), .B2(new_n762_), .ZN(G1332gat));
  OAI21_X1  g562(.A(G64gat), .B1(new_n749_), .B2(new_n471_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT48), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n471_), .A2(G64gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n759_), .B2(new_n766_), .ZN(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n749_), .B2(new_n688_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT49), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n688_), .A2(G71gat), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT111), .Z(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n759_), .B2(new_n771_), .ZN(G1334gat));
  OAI21_X1  g571(.A(G78gat), .B1(new_n749_), .B2(new_n447_), .ZN(new_n773_));
  XOR2_X1   g572(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n447_), .A2(G78gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n759_), .B2(new_n776_), .ZN(G1335gat));
  NOR3_X1   g576(.A1(new_n754_), .A2(new_n646_), .A3(new_n599_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n713_), .A2(KEYINPUT113), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n713_), .A2(KEYINPUT113), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n530_), .B1(new_n782_), .B2(new_n639_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n699_), .A2(new_n754_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n757_), .A2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(G85gat), .A3(new_n396_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT114), .B1(new_n783_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788_));
  INV_X1    g587(.A(new_n786_), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n396_), .B(new_n779_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n788_), .B(new_n789_), .C1(new_n790_), .C2(new_n530_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(G1336gat));
  INV_X1    g591(.A(new_n785_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n531_), .A3(new_n659_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n782_), .A2(new_n659_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n531_), .ZN(G1337gat));
  INV_X1    g595(.A(G99gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n782_), .B2(new_n259_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(new_n259_), .A3(new_n520_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT51), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n688_), .B(new_n779_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n802_), .B(new_n799_), .C1(new_n803_), .C2(new_n797_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n793_), .A2(new_n451_), .A3(new_n521_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n778_), .A2(new_n451_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n476_), .A2(KEYINPUT43), .A3(new_n704_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n711_), .B1(new_n710_), .B2(new_n703_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT115), .B(new_n808_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G106gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n807_), .B1(new_n705_), .B2(new_n712_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT115), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n812_), .A2(new_n814_), .A3(KEYINPUT52), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n713_), .A2(new_n808_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G106gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n813_), .B2(KEYINPUT115), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n816_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n806_), .B1(new_n815_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT53), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n806_), .C1(new_n815_), .C2(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1339gat));
  NAND3_X1  g626(.A1(new_n473_), .A2(new_n259_), .A3(new_n639_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n617_), .B1(new_n550_), .B2(new_n612_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n608_), .A2(KEYINPUT117), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n830_), .A2(KEYINPUT55), .A3(new_n605_), .A4(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(new_n626_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(KEYINPUT55), .A3(new_n605_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n614_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n835_), .B(new_n831_), .C1(new_n836_), .C2(KEYINPUT55), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n834_), .A2(new_n837_), .A3(KEYINPUT56), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n837_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n519_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n840_));
  OAI22_X1  g639(.A1(new_n838_), .A2(new_n839_), .B1(new_n840_), .B2(KEYINPUT116), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n629_), .A2(new_n646_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n829_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n834_), .A2(new_n837_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n834_), .A2(new_n837_), .A3(KEYINPUT56), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n843_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n840_), .A2(KEYINPUT116), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(KEYINPUT118), .A4(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n514_), .A2(G229gat), .A3(G233gat), .A4(new_n493_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n505_), .A2(new_n493_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n509_), .B1(new_n855_), .B2(new_n494_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n511_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n631_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n845_), .A2(new_n853_), .A3(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(KEYINPUT57), .A3(new_n643_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n850_), .A2(new_n629_), .A3(new_n857_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n862_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n703_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n859_), .B2(new_n643_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n860_), .B(new_n865_), .C1(new_n866_), .C2(KEYINPUT119), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n868_), .A2(new_n829_), .B1(new_n631_), .B2(new_n857_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n644_), .B1(new_n869_), .B2(new_n853_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n870_), .A2(new_n871_), .A3(KEYINPUT57), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n598_), .B1(new_n867_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n636_), .B2(new_n519_), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n601_), .A2(KEYINPUT54), .A3(new_n646_), .A4(new_n635_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n828_), .B1(new_n873_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(G113gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n646_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n828_), .A2(KEYINPUT59), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n860_), .A2(new_n865_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n598_), .B1(new_n883_), .B2(new_n866_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n884_), .A2(KEYINPUT121), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n877_), .B1(new_n884_), .B2(KEYINPUT121), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n879_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n871_), .B1(new_n870_), .B2(KEYINPUT57), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n866_), .A2(KEYINPUT119), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n860_), .A4(new_n865_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n877_), .B1(new_n893_), .B2(new_n598_), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n894_), .C2(new_n828_), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n519_), .B(new_n887_), .C1(new_n890_), .C2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n881_), .B1(new_n896_), .B2(new_n880_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n754_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n879_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n754_), .B(new_n887_), .C1(new_n890_), .C2(new_n895_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n898_), .ZN(G1341gat));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n879_), .A2(new_n903_), .A3(new_n599_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n598_), .B(new_n887_), .C1(new_n890_), .C2(new_n895_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1342gat));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n879_), .A2(new_n907_), .A3(new_n644_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n704_), .B(new_n887_), .C1(new_n890_), .C2(new_n895_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1343gat));
  NOR2_X1   g709(.A1(new_n894_), .A2(new_n447_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n659_), .A2(new_n259_), .A3(new_n396_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n646_), .A3(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n635_), .A3(new_n912_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n911_), .A2(new_n917_), .A3(new_n599_), .A4(new_n912_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n873_), .A2(new_n878_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n919_), .A2(new_n451_), .A3(new_n599_), .A4(new_n912_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT122), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n921_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1346gat));
  NAND2_X1  g723(.A1(new_n911_), .A2(new_n912_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G162gat), .B1(new_n925_), .B2(new_n704_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n643_), .A2(G162gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(G1347gat));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n885_), .A2(new_n886_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n475_), .A2(new_n659_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n451_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n519_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n929_), .B1(new_n934_), .B2(new_n219_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n241_), .ZN(new_n936_));
  OAI211_X1 g735(.A(KEYINPUT62), .B(G169gat), .C1(new_n933_), .C2(new_n519_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(G1348gat));
  INV_X1    g737(.A(new_n933_), .ZN(new_n939_));
  AOI21_X1  g738(.A(G176gat), .B1(new_n939_), .B2(new_n635_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n451_), .B1(new_n873_), .B2(new_n878_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n931_), .A2(new_n220_), .A3(new_n754_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1349gat));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n475_), .A2(new_n659_), .A3(new_n599_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n919_), .A2(new_n447_), .A3(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n941_), .A2(KEYINPUT123), .A3(new_n946_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n206_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n210_), .A2(new_n362_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n599_), .A2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n933_), .A2(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n944_), .B1(new_n951_), .B2(new_n954_), .ZN(new_n955_));
  NOR4_X1   g754(.A1(new_n894_), .A2(new_n948_), .A3(new_n451_), .A4(new_n945_), .ZN(new_n956_));
  AOI21_X1  g755(.A(KEYINPUT123), .B1(new_n941_), .B2(new_n946_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n232_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n933_), .A2(new_n953_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n958_), .A2(new_n959_), .A3(KEYINPUT124), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n955_), .A2(new_n960_), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n933_), .B2(new_n704_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n644_), .A2(new_n209_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n962_), .B1(new_n933_), .B2(new_n963_), .ZN(G1351gat));
  NOR3_X1   g763(.A1(new_n471_), .A2(new_n259_), .A3(new_n639_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n911_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n966_), .A2(new_n519_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(new_n317_), .ZN(G1352gat));
  NOR2_X1   g767(.A1(new_n966_), .A2(new_n754_), .ZN(new_n969_));
  XOR2_X1   g768(.A(KEYINPUT125), .B(G204gat), .Z(new_n970_));
  XNOR2_X1  g769(.A(new_n969_), .B(new_n970_), .ZN(G1353gat));
  INV_X1    g770(.A(new_n966_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n598_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n975_), .B(KEYINPUT126), .ZN(new_n976_));
  INV_X1    g775(.A(new_n976_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n974_), .A2(new_n977_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n972_), .A2(new_n976_), .A3(new_n973_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n966_), .B2(new_n704_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n644_), .A2(new_n311_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n966_), .B2(new_n982_), .ZN(G1355gat));
endmodule


