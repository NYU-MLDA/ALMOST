//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT92), .ZN(new_n203_));
  XOR2_X1   g002(.A(G197gat), .B(G204gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT21), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n203_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT3), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(KEYINPUT1), .B2(new_n220_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(KEYINPUT1), .B2(new_n220_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n217_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(new_n215_), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n219_), .A2(new_n223_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n212_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G78gat), .ZN(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(G78gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n233_), .B(new_n212_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n214_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n214_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n235_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G22gat), .B(G50gat), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n228_), .A2(new_n229_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n246_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n244_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT93), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n250_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n242_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n238_), .A2(new_n241_), .A3(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  AND3_X1   g059(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n263_), .A2(new_n264_), .B1(G169gat), .B2(G176gat), .ZN(new_n265_));
  INV_X1    g064(.A(G176gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT87), .ZN(new_n267_));
  INV_X1    g066(.A(G169gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT22), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT22), .B(G169gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n266_), .B(new_n269_), .C1(new_n270_), .C2(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n273_), .A2(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT24), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(new_n268_), .A3(new_n266_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n272_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n260_), .B1(new_n288_), .B2(new_n212_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT19), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT96), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n270_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n266_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n265_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT95), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT94), .B1(new_n263_), .B2(new_n280_), .ZN(new_n299_));
  AND4_X1   g098(.A1(KEYINPUT94), .A2(new_n280_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n298_), .B(new_n278_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT94), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n285_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n263_), .A2(KEYINPUT94), .A3(new_n280_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n298_), .B1(new_n306_), .B2(new_n278_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n297_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n308_), .A2(KEYINPUT98), .A3(new_n212_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT98), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n263_), .A2(new_n264_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n277_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n295_), .B2(new_n266_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n278_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT95), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n315_), .B2(new_n301_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n210_), .A2(new_n211_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n310_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n293_), .B1(new_n309_), .B2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n212_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n308_), .B2(new_n212_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT97), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n292_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n272_), .A2(new_n287_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n260_), .B1(new_n324_), .B2(new_n317_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT97), .B1(new_n326_), .B2(new_n291_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n319_), .B1(new_n323_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n332_), .B(new_n319_), .C1(new_n323_), .C2(new_n327_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT99), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT99), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n328_), .A2(new_n338_), .A3(new_n333_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n297_), .A2(new_n317_), .A3(new_n314_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n292_), .B1(new_n341_), .B2(new_n289_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n321_), .B2(new_n292_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n335_), .B(KEYINPUT27), .C1(new_n332_), .C2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT104), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G57gat), .B(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT100), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G134gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n221_), .B(new_n222_), .C1(new_n216_), .C2(new_n218_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n225_), .A2(new_n227_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n354_), .B(new_n355_), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n228_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n361_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n228_), .A2(new_n360_), .A3(KEYINPUT4), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n353_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n352_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n350_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n364_), .A2(new_n350_), .A3(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n345_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(KEYINPUT104), .A3(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(G71gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G99gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n288_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(new_n360_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G15gat), .B(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT88), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT30), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT31), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n378_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n372_), .A2(new_n384_), .ZN(new_n385_));
  AND4_X1   g184(.A1(new_n259_), .A2(new_n340_), .A3(new_n344_), .A4(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n387_));
  NAND3_X1  g186(.A1(new_n362_), .A2(new_n363_), .A3(new_n353_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n359_), .A2(new_n361_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n350_), .B1(new_n389_), .B2(new_n352_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n366_), .A2(new_n387_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT33), .B(new_n350_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT102), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n393_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n391_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n328_), .B1(KEYINPUT32), .B2(new_n332_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n399_));
  OAI22_X1  g198(.A1(new_n367_), .A2(new_n368_), .B1(new_n399_), .B2(new_n343_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n259_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n259_), .A2(new_n372_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n340_), .A2(new_n403_), .A3(new_n344_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n383_), .B(KEYINPUT89), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n386_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G1gat), .A2(G8gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G1gat), .A2(G8gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT79), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(G1gat), .A2(G8gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G15gat), .ZN(new_n417_));
  INV_X1    g216(.A(G22gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G15gat), .A2(G22gat), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n419_), .A2(new_n420_), .B1(KEYINPUT14), .B2(new_n409_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n424_));
  INV_X1    g223(.A(G36gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G29gat), .ZN(new_n426_));
  INV_X1    g225(.A(G29gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G36gat), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n426_), .A2(new_n428_), .A3(KEYINPUT73), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT73), .B1(new_n426_), .B2(new_n428_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G43gat), .B(G50gat), .Z(new_n431_));
  NOR3_X1   g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G43gat), .B(G50gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT73), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n427_), .A2(G36gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n425_), .A2(G29gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n426_), .A2(new_n428_), .A3(KEYINPUT73), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n433_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n423_), .B(new_n424_), .C1(new_n432_), .C2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n438_), .A3(new_n433_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n431_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n421_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n419_), .A2(new_n420_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n409_), .A2(KEYINPUT14), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n412_), .A2(new_n415_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n441_), .B(new_n442_), .C1(new_n443_), .C2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n440_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G229gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n440_), .A2(new_n447_), .A3(KEYINPUT83), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n442_), .A2(new_n441_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT15), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n442_), .A2(new_n441_), .A3(KEYINPUT15), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n457_), .B(new_n458_), .C1(new_n443_), .C2(new_n446_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n451_), .A3(new_n440_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G113gat), .B(G141gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT84), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G169gat), .B(G197gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n454_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n467_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n454_), .A2(new_n460_), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n468_), .A2(new_n469_), .B1(new_n470_), .B2(new_n464_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n466_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT86), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n470_), .A2(new_n464_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n408_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G190gat), .B(G218gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G134gat), .B(G162gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT65), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n487_));
  AND2_X1   g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT10), .B(G99gat), .ZN(new_n491_));
  OAI22_X1  g290(.A1(new_n489_), .A2(new_n490_), .B1(G106gat), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT64), .ZN(new_n493_));
  OAI211_X1 g292(.A(G85gat), .B(G92gat), .C1(new_n493_), .C2(KEYINPUT9), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n493_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n493_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G99gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n232_), .A3(KEYINPUT7), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(G99gat), .B2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n506_));
  AND2_X1   g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n505_), .A2(new_n506_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n506_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n499_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n458_), .A3(new_n457_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n516_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n455_), .B(new_n499_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT75), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n520_), .A2(new_n517_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT74), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n522_), .A2(new_n529_), .A3(new_n523_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n516_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n527_), .B(new_n528_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n524_), .A2(KEYINPUT74), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(new_n530_), .A3(new_n516_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n527_), .B1(new_n536_), .B2(new_n528_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n483_), .B(new_n526_), .C1(new_n534_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n482_), .B(KEYINPUT36), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n526_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(KEYINPUT78), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n528_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT75), .ZN(new_n545_));
  AOI211_X1 g344(.A(KEYINPUT78), .B(new_n525_), .C1(new_n545_), .C2(new_n533_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n539_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n538_), .A2(KEYINPUT76), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT77), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n550_), .A3(new_n540_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n525_), .B1(new_n545_), .B2(new_n533_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT76), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n483_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n541_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT37), .B1(new_n556_), .B2(new_n550_), .ZN(new_n557_));
  OAI22_X1  g356(.A1(new_n548_), .A2(KEYINPUT37), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n560_));
  NOR2_X1   g359(.A1(new_n492_), .A2(new_n498_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n506_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n484_), .A2(KEYINPUT65), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n566_), .A2(new_n567_), .B1(new_n503_), .B2(new_n501_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n562_), .B1(new_n568_), .B2(new_n511_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n505_), .A2(new_n506_), .A3(new_n512_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n561_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G57gat), .B(G64gat), .Z(new_n572_));
  INV_X1    g371(.A(KEYINPUT11), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT67), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n573_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G71gat), .B(G78gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT67), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT11), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .A4(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n576_), .B1(KEYINPUT11), .B2(new_n577_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT11), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n578_), .B1(new_n577_), .B2(KEYINPUT11), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n581_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n560_), .B1(new_n571_), .B2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n580_), .A2(new_n584_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n515_), .A2(KEYINPUT12), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n585_), .B(new_n499_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n589_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n590_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n571_), .A2(new_n585_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT5), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT69), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(KEYINPUT70), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT71), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT70), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n606_), .A3(new_n601_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n605_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n559_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT71), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(KEYINPUT13), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n585_), .B(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n443_), .A2(new_n446_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT82), .ZN(new_n623_));
  XOR2_X1   g422(.A(G127gat), .B(G155gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT17), .Z(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n622_), .A2(KEYINPUT81), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT81), .B1(new_n622_), .B2(new_n631_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n630_), .A2(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n558_), .A2(new_n616_), .A3(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n479_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n372_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(G1gat), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT38), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n408_), .A2(new_n548_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n635_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT106), .B1(new_n615_), .B2(new_n477_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n648_), .B(new_n478_), .C1(new_n610_), .C2(new_n614_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n645_), .A2(new_n646_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n372_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n644_), .B1(new_n652_), .B2(G1gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n643_), .B1(new_n653_), .B2(new_n640_), .ZN(G1324gat));
  NAND2_X1  g453(.A1(new_n340_), .A2(new_n344_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n645_), .A2(new_n655_), .A3(new_n646_), .A4(new_n650_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT107), .B1(new_n656_), .B2(G8gat), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  INV_X1    g460(.A(G8gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n637_), .A2(new_n662_), .A3(new_n655_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .A4(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n664_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n661_), .A2(new_n663_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n669_), .ZN(G1325gat));
  AOI21_X1  g469(.A(new_n417_), .B1(new_n651_), .B2(new_n406_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT41), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n637_), .A2(new_n417_), .A3(new_n406_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(new_n259_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n418_), .B1(new_n651_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT42), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n637_), .A2(new_n418_), .A3(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n548_), .A2(new_n635_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n616_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n479_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G29gat), .B1(new_n683_), .B2(new_n372_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n558_), .B2(KEYINPUT109), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n549_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT37), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n542_), .A2(new_n540_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(KEYINPUT77), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT78), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n540_), .B1(new_n552_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n538_), .B1(new_n692_), .B2(new_n546_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n687_), .A2(new_n690_), .B1(new_n693_), .B2(new_n688_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n686_), .B1(new_n408_), .B2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n406_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n696_));
  OAI221_X1 g495(.A(new_n558_), .B1(KEYINPUT109), .B2(new_n685_), .C1(new_n696_), .C2(new_n386_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n608_), .A2(new_n609_), .A3(new_n559_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT13), .B1(new_n612_), .B2(new_n613_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n477_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n648_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n615_), .A2(KEYINPUT106), .A3(new_n477_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n635_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n698_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n707_), .B(new_n704_), .C1(new_n695_), .C2(new_n697_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n638_), .A2(new_n427_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n684_), .B1(new_n709_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n425_), .B1(new_n709_), .B2(new_n655_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n655_), .A2(new_n425_), .ZN(new_n715_));
  OR3_X1    g514(.A1(new_n682_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n682_), .B2(new_n715_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n712_), .B1(new_n713_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n718_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n655_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n706_), .A2(new_n708_), .A3(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n720_), .B(KEYINPUT46), .C1(new_n722_), .C2(new_n425_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n719_), .A2(new_n723_), .ZN(G1329gat));
  INV_X1    g523(.A(new_n706_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n698_), .A2(new_n705_), .A3(KEYINPUT44), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n383_), .A2(G43gat), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G43gat), .B1(new_n683_), .B2(new_n406_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT47), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n709_), .B2(new_n727_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1330gat));
  OR3_X1    g533(.A1(new_n682_), .A2(G50gat), .A3(new_n259_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n675_), .A3(new_n726_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT111), .B1(new_n736_), .B2(G50gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n408_), .A2(new_n615_), .A3(new_n477_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n558_), .A2(new_n635_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n372_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n615_), .A2(new_n635_), .A3(new_n477_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n645_), .A2(G57gat), .A3(new_n372_), .A4(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n746_), .A2(new_n747_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n744_), .A2(new_n748_), .A3(new_n749_), .ZN(G1332gat));
  NAND2_X1  g549(.A1(new_n645_), .A2(new_n745_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G64gat), .B1(new_n751_), .B2(new_n721_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n721_), .A2(G64gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n742_), .B2(new_n755_), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n751_), .B2(new_n407_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT49), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n743_), .A2(new_n374_), .A3(new_n406_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1334gat));
  OAI21_X1  g559(.A(G78gat), .B1(new_n751_), .B2(new_n259_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT50), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n675_), .A2(new_n233_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT114), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n742_), .B2(new_n764_), .ZN(G1335gat));
  INV_X1    g564(.A(G85gat), .ZN(new_n766_));
  INV_X1    g565(.A(new_n680_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n740_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n768_), .B2(new_n638_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT115), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n616_), .A2(new_n635_), .A3(new_n478_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n638_), .A2(new_n766_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(G1336gat));
  INV_X1    g573(.A(new_n768_), .ZN(new_n775_));
  INV_X1    g574(.A(G92gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n655_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n772_), .A2(new_n655_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n776_), .ZN(G1337gat));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n384_), .A2(new_n491_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT116), .B1(new_n768_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n772_), .A2(new_n406_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n788_), .A2(new_n500_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n789_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n786_), .A3(new_n792_), .A4(new_n785_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n775_), .A2(new_n232_), .A3(new_n675_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n772_), .A2(new_n675_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G106gat), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT52), .B(new_n232_), .C1(new_n772_), .C2(new_n675_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n795_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  INV_X1    g603(.A(G113gat), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n690_), .A2(new_n551_), .A3(new_n549_), .A4(new_n554_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n693_), .A2(new_n688_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n635_), .A2(new_n477_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n806_), .A2(new_n615_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n810_));
  NOR2_X1   g609(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n694_), .A2(new_n615_), .A3(new_n808_), .A4(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n451_), .B1(new_n619_), .B2(new_n455_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n464_), .B1(new_n459_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n612_), .A2(new_n613_), .A3(new_n465_), .A4(new_n819_), .ZN(new_n820_));
  AND4_X1   g619(.A1(new_n589_), .A2(new_n586_), .A3(new_n588_), .A4(new_n590_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n586_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n592_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(KEYINPUT55), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n822_), .A2(new_n825_), .A3(new_n592_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n601_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT56), .B(new_n601_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n829_), .A2(KEYINPUT119), .A3(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n477_), .B(new_n603_), .C1(KEYINPUT119), .C2(new_n830_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n820_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n693_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n603_), .A2(new_n465_), .A3(new_n819_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n830_), .A2(KEYINPUT120), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n829_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n830_), .A2(KEYINPUT120), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT58), .B(new_n837_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n558_), .A3(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n833_), .A2(KEYINPUT57), .A3(new_n693_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n836_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n815_), .B1(new_n847_), .B2(new_n635_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n655_), .A2(new_n675_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n372_), .A3(new_n383_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n805_), .B1(new_n853_), .B2(new_n478_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT121), .B(new_n805_), .C1(new_n853_), .C2(new_n478_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n829_), .A2(KEYINPUT119), .A3(new_n830_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n830_), .A2(KEYINPUT119), .ZN(new_n861_));
  INV_X1    g660(.A(new_n603_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n864_));
  AOI211_X1 g663(.A(new_n835_), .B(new_n548_), .C1(new_n864_), .C2(new_n820_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n833_), .B2(new_n693_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n646_), .B1(new_n867_), .B2(new_n845_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT59), .B(new_n852_), .C1(new_n868_), .C2(new_n815_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n859_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n478_), .A2(new_n805_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n856_), .A2(new_n857_), .B1(new_n870_), .B2(new_n871_), .ZN(G1340gat));
  NOR2_X1   g671(.A1(new_n615_), .A2(KEYINPUT60), .ZN(new_n873_));
  MUX2_X1   g672(.A(new_n873_), .B(KEYINPUT60), .S(G120gat), .Z(new_n874_));
  NAND3_X1  g673(.A1(new_n849_), .A2(new_n852_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n615_), .B1(new_n859_), .B2(new_n869_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G120gat), .B1(new_n876_), .B2(KEYINPUT122), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n878_), .B(new_n615_), .C1(new_n859_), .C2(new_n869_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n877_), .B2(new_n879_), .ZN(G1341gat));
  AOI21_X1  g679(.A(new_n635_), .B1(new_n859_), .B2(new_n869_), .ZN(new_n881_));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n646_), .A2(new_n882_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n881_), .A2(new_n882_), .B1(new_n853_), .B2(new_n883_), .ZN(G1342gat));
  AOI21_X1  g683(.A(new_n694_), .B1(new_n859_), .B2(new_n869_), .ZN(new_n885_));
  INV_X1    g684(.A(G134gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n548_), .A2(new_n886_), .ZN(new_n887_));
  OAI22_X1  g686(.A1(new_n885_), .A2(new_n886_), .B1(new_n853_), .B2(new_n887_), .ZN(G1343gat));
  NAND4_X1  g687(.A1(new_n721_), .A2(new_n407_), .A3(new_n372_), .A4(new_n675_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT123), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n849_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n477_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n616_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g694(.A1(new_n849_), .A2(new_n890_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n635_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT61), .B(G155gat), .Z(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n896_), .B2(new_n694_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n693_), .A2(G162gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n896_), .B2(new_n901_), .ZN(G1347gat));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903_));
  NOR4_X1   g702(.A1(new_n721_), .A2(new_n407_), .A3(new_n372_), .A4(new_n675_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n477_), .B(new_n904_), .C1(new_n868_), .C2(new_n815_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n849_), .A2(new_n295_), .A3(new_n477_), .A4(new_n904_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT62), .B1(new_n905_), .B2(G169gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n903_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(G169gat), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n913_), .A2(KEYINPUT124), .A3(new_n907_), .A4(new_n906_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(G1348gat));
  INV_X1    g714(.A(new_n904_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n848_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n616_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n646_), .ZN(new_n920_));
  MUX2_X1   g719(.A(new_n273_), .B(G183gat), .S(new_n920_), .Z(G1350gat));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n274_), .A3(new_n548_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n848_), .A2(new_n694_), .A3(new_n916_), .ZN(new_n923_));
  INV_X1    g722(.A(G190gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n407_), .A2(new_n403_), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT125), .Z(new_n927_));
  NOR3_X1   g726(.A1(new_n848_), .A2(new_n721_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n477_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n616_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g731(.A(new_n635_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n928_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT126), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT127), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n934_), .B(new_n937_), .ZN(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n928_), .A2(new_n939_), .A3(new_n548_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n928_), .A2(new_n558_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n939_), .ZN(G1355gat));
endmodule


