//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(G15gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT30), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT80), .B(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT79), .ZN(new_n208_));
  INV_X1    g007(.A(G169gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT22), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(KEYINPUT22), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n207_), .B(new_n210_), .C1(new_n211_), .C2(new_n208_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT23), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(KEYINPUT82), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n218_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n224_), .B(KEYINPUT23), .C1(new_n217_), .C2(new_n218_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT81), .B1(new_n212_), .B2(new_n213_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n216_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT78), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT78), .B1(new_n217_), .B2(KEYINPUT25), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n234_));
  OR2_X1    g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  MUX2_X1   g034(.A(KEYINPUT24), .B(new_n234_), .S(new_n235_), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n219_), .A2(new_n221_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT83), .B1(new_n228_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n227_), .A2(new_n226_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n215_), .B2(new_n214_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n239_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247_));
  INV_X1    g046(.A(G43gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G113gat), .B(G120gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n246_), .A2(new_n249_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n206_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n256_), .A3(new_n205_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G78gat), .B(G106gat), .ZN(new_n263_));
  INV_X1    g062(.A(G228gat), .ZN(new_n264_));
  INV_X1    g063(.A(G233gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G197gat), .B(G204gat), .Z(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT21), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT21), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n271_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT84), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT85), .B1(new_n276_), .B2(KEYINPUT1), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT84), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n275_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT85), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n276_), .A2(KEYINPUT1), .ZN(new_n283_));
  OR2_X1    g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n277_), .A2(new_n282_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G141gat), .B(G148gat), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OR3_X1    g086(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289_));
  INV_X1    g088(.A(G141gat), .ZN(new_n290_));
  INV_X1    g089(.A(G148gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n288_), .A2(new_n292_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(new_n276_), .A3(new_n284_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n287_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT86), .ZN(new_n298_));
  INV_X1    g097(.A(new_n296_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT86), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n267_), .B(new_n274_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n267_), .B1(new_n306_), .B2(new_n274_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT88), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n274_), .A2(new_n267_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n300_), .A2(new_n301_), .ZN(new_n311_));
  AOI211_X1 g110(.A(KEYINPUT86), .B(new_n299_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n313_), .B2(KEYINPUT29), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n307_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n263_), .B1(new_n309_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n305_), .A2(new_n308_), .A3(KEYINPUT88), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n315_), .B1(new_n314_), .B2(new_n307_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n263_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(KEYINPUT87), .A3(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT28), .B1(new_n313_), .B2(KEYINPUT29), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n303_), .A2(new_n324_), .A3(new_n304_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G22gat), .B(G50gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n322_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n318_), .A2(new_n319_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n263_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n330_), .B1(new_n335_), .B2(new_n321_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n262_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n322_), .A2(new_n331_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n259_), .A2(new_n261_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n321_), .A3(new_n330_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n274_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n229_), .A2(new_n232_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n236_), .A2(new_n225_), .A3(new_n222_), .A4(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n207_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n213_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(KEYINPUT89), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n237_), .A2(new_n223_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n352_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n346_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT20), .B1(new_n355_), .B2(new_n274_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n344_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n240_), .A2(new_n245_), .A3(new_n343_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n355_), .B2(new_n274_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n360_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT18), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n359_), .B1(new_n344_), .B2(new_n356_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n370_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT98), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT98), .ZN(new_n377_));
  AOI211_X1 g176(.A(new_n377_), .B(new_n370_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT27), .B(new_n371_), .C1(new_n376_), .C2(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n344_), .A2(new_n359_), .A3(new_n356_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n375_), .B1(new_n380_), .B2(new_n365_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n371_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G57gat), .B(G85gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT94), .ZN(new_n387_));
  XOR2_X1   g186(.A(G1gat), .B(G29gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT92), .B(KEYINPUT4), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n313_), .A2(new_n253_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT91), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n298_), .A2(new_n398_), .A3(new_n302_), .A4(new_n253_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n311_), .A2(new_n312_), .A3(new_n254_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT90), .B1(new_n297_), .B2(new_n253_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n397_), .B1(new_n402_), .B2(KEYINPUT4), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n395_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n392_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT97), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n402_), .A2(KEYINPUT4), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n404_), .B(new_n391_), .C1(new_n408_), .C2(new_n397_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n407_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n385_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n382_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT95), .B1(new_n409_), .B2(new_n413_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n404_), .A2(new_n391_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n403_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT33), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n394_), .A2(new_n395_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT96), .B1(new_n408_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n402_), .A2(KEYINPUT4), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT96), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n391_), .B1(new_n402_), .B2(new_n396_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n414_), .A2(new_n415_), .A3(new_n419_), .A4(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n374_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n380_), .A2(new_n365_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n391_), .B1(new_n432_), .B2(new_n404_), .ZN(new_n433_));
  OAI221_X1 g232(.A(new_n429_), .B1(new_n431_), .B2(new_n428_), .C1(new_n433_), .C2(new_n417_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n338_), .A2(new_n262_), .A3(new_n340_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n342_), .A2(new_n412_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G232gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT34), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT35), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G29gat), .B(G36gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT68), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G43gat), .B(G50gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n444_), .A2(KEYINPUT68), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(KEYINPUT68), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n446_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT15), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT10), .B(G99gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT64), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G85gat), .A2(G92gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI221_X1 g268(.A(new_n459_), .B1(G106gat), .B2(new_n460_), .C1(new_n463_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n457_), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT65), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n456_), .A2(new_n458_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n474_), .A2(new_n476_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n466_), .A2(new_n468_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n471_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  AOI211_X1 g285(.A(KEYINPUT8), .B(new_n484_), .C1(new_n482_), .C2(new_n459_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n470_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n454_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n448_), .A2(new_n451_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT66), .B(new_n470_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n441_), .A2(new_n442_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n443_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n489_), .B(KEYINPUT69), .ZN(new_n500_));
  INV_X1    g299(.A(new_n443_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G190gat), .B(G218gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT36), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n505_), .B(KEYINPUT36), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n438_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G57gat), .B(G64gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT11), .ZN(new_n515_));
  XOR2_X1   g314(.A(G71gat), .B(G78gat), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n514_), .A2(KEYINPUT11), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n515_), .A2(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(G231gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT70), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G1gat), .A2(G8gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT14), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G8gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT74), .ZN(new_n533_));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT17), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n524_), .B(new_n530_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n532_), .A2(KEYINPUT71), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n533_), .A2(new_n539_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n521_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n488_), .A2(new_n548_), .A3(KEYINPUT12), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n521_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(KEYINPUT12), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n493_), .A2(new_n495_), .A3(new_n521_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT67), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n551_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n482_), .A2(new_n459_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n471_), .A3(new_n485_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n480_), .A2(new_n481_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(KEYINPUT65), .B2(new_n459_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n484_), .B1(new_n562_), .B2(new_n476_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n560_), .B1(new_n563_), .B2(new_n471_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT66), .B1(new_n564_), .B2(new_n470_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n495_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n548_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n553_), .B1(new_n567_), .B2(new_n552_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n558_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT5), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n558_), .B2(new_n568_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(KEYINPUT13), .A3(new_n576_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n530_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n494_), .A2(KEYINPUT75), .A3(new_n530_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n494_), .B2(new_n530_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n452_), .A2(new_n453_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT15), .B1(new_n448_), .B2(new_n451_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n531_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT76), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n586_), .A2(new_n593_), .A3(new_n594_), .A4(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n586_), .A2(new_n593_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n594_), .B1(new_n597_), .B2(new_n588_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT77), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT77), .B(new_n602_), .C1(new_n596_), .C2(new_n598_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n581_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n513_), .A2(new_n547_), .A3(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n410_), .A2(new_n411_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT99), .Z(new_n613_));
  NOR3_X1   g412(.A1(new_n332_), .A2(new_n336_), .A3(new_n262_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n339_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n412_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n435_), .A2(new_n437_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n511_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n507_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT37), .B1(new_n508_), .B2(new_n511_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n533_), .A2(new_n539_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n545_), .A2(new_n546_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n618_), .A2(new_n609_), .A3(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n628_), .A2(G1gat), .A3(new_n611_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT38), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n613_), .A2(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(new_n385_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G8gat), .B1(new_n610_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT39), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n632_), .A2(G8gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n628_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  OAI21_X1  g437(.A(G15gat), .B1(new_n610_), .B2(new_n262_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT100), .Z(new_n640_));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n628_), .A2(G15gat), .A3(new_n262_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT101), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n642_), .A2(new_n643_), .A3(new_n645_), .ZN(G1326gat));
  NOR2_X1   g445(.A1(new_n332_), .A2(new_n336_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G22gat), .B1(new_n610_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n647_), .A2(G22gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n628_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1327gat));
  INV_X1    g452(.A(new_n512_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n547_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT97), .B1(new_n433_), .B2(new_n417_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n406_), .A2(new_n409_), .A3(new_n407_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n384_), .A4(new_n379_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n436_), .B1(new_n427_), .B2(new_n434_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n609_), .B(new_n655_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n618_), .A2(KEYINPUT104), .A3(new_n609_), .A4(new_n655_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n611_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n623_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT103), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n618_), .A2(new_n671_), .A3(new_n668_), .A4(new_n623_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n621_), .A2(new_n622_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n438_), .B2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n608_), .A2(new_n547_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n676_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n666_), .A2(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n667_), .B1(new_n681_), .B2(new_n682_), .ZN(G1328gat));
  NOR2_X1   g482(.A1(new_n632_), .A2(G36gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n663_), .A2(new_n664_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n688_));
  NAND4_X1  g487(.A1(new_n663_), .A2(new_n664_), .A3(KEYINPUT106), .A4(new_n684_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n679_), .A2(new_n385_), .A3(new_n680_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G36gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n692_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1329gat));
  NOR2_X1   g497(.A1(new_n262_), .A2(new_n248_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n679_), .A2(new_n680_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT108), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n679_), .A2(new_n702_), .A3(new_n680_), .A4(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n665_), .A2(new_n339_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT109), .B(G43gat), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(new_n703_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n701_), .A2(new_n709_), .A3(new_n703_), .A4(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1330gat));
  INV_X1    g510(.A(new_n647_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G50gat), .B1(new_n665_), .B2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n681_), .B2(new_n714_), .ZN(G1331gat));
  NAND2_X1  g514(.A1(new_n547_), .A2(new_n673_), .ZN(new_n716_));
  NOR4_X1   g515(.A1(new_n438_), .A2(new_n607_), .A3(new_n581_), .A4(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n666_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n626_), .A2(new_n581_), .A3(new_n607_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n513_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n611_), .A2(KEYINPUT110), .ZN(new_n722_));
  MUX2_X1   g521(.A(KEYINPUT110), .B(new_n722_), .S(G57gat), .Z(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n721_), .B2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g523(.A(G64gat), .B1(new_n720_), .B2(new_n632_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n717_), .A2(new_n728_), .A3(new_n385_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n720_), .B2(new_n262_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT49), .ZN(new_n733_));
  INV_X1    g532(.A(G71gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n717_), .A2(new_n734_), .A3(new_n339_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n720_), .B2(new_n647_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT50), .ZN(new_n738_));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n717_), .A2(new_n739_), .A3(new_n712_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n438_), .A2(new_n607_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n581_), .A2(new_n547_), .A3(new_n654_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n464_), .B1(new_n744_), .B2(new_n611_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT113), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n581_), .A2(new_n547_), .A3(new_n607_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n675_), .A2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n611_), .A2(new_n464_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(G1336gat));
  INV_X1    g549(.A(new_n744_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n465_), .A3(new_n385_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n748_), .A2(new_n385_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n465_), .ZN(G1337gat));
  OR3_X1    g553(.A1(new_n744_), .A2(new_n460_), .A3(new_n262_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n748_), .A2(new_n339_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT114), .B(new_n755_), .C1(new_n756_), .C2(new_n478_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g557(.A1(new_n751_), .A2(new_n479_), .A3(new_n712_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n675_), .A2(new_n712_), .A3(new_n747_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G106gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G106gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g564(.A1(new_n586_), .A2(new_n593_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT76), .B1(new_n766_), .B2(new_n589_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(new_n590_), .A3(new_n595_), .A4(new_n602_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n587_), .A2(new_n588_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT118), .B1(new_n769_), .B2(new_n603_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n584_), .A2(new_n585_), .B1(new_n452_), .B2(new_n531_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT118), .B(new_n603_), .C1(new_n771_), .C2(new_n589_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n588_), .B2(new_n766_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n569_), .B2(new_n574_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  INV_X1    g575(.A(new_n549_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT12), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n567_), .B2(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n552_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n556_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  INV_X1    g582(.A(new_n553_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n552_), .B(new_n549_), .C1(new_n550_), .C2(KEYINPUT12), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n782_), .A2(new_n783_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n779_), .B(KEYINPUT55), .C1(new_n780_), .C2(new_n781_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n776_), .B(new_n574_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n782_), .A2(new_n783_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n784_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n787_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n573_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n775_), .B1(new_n788_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n775_), .B(KEYINPUT58), .C1(new_n788_), .C2(new_n792_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n623_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n606_), .B1(new_n569_), .B2(new_n574_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT117), .B1(new_n776_), .B2(KEYINPUT116), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n790_), .B1(new_n558_), .B2(KEYINPUT55), .ZN(new_n800_));
  INV_X1    g599(.A(new_n787_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n573_), .B(new_n799_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n574_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n776_), .A2(KEYINPUT116), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n803_), .B2(KEYINPUT56), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n798_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n774_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n512_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n797_), .B1(new_n811_), .B2(KEYINPUT57), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n813_), .B(new_n512_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n626_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n627_), .A2(new_n606_), .A3(new_n581_), .A4(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n581_), .A2(new_n606_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n716_), .B2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n611_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n341_), .A2(new_n385_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n607_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n815_), .A2(new_n821_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n666_), .A4(new_n823_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n822_), .A2(new_n827_), .A3(KEYINPUT59), .A4(new_n823_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n607_), .A2(G113gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n825_), .B1(new_n835_), .B2(new_n836_), .ZN(G1340gat));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n581_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n824_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n581_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n838_), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n824_), .B2(new_n547_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n547_), .A2(G127gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n835_), .B2(new_n844_), .ZN(G1342gat));
  AOI21_X1  g644(.A(G134gat), .B1(new_n824_), .B2(new_n512_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n623_), .A2(G134gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n835_), .B2(new_n847_), .ZN(G1343gat));
  NAND3_X1  g647(.A1(new_n822_), .A2(new_n615_), .A3(new_n632_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n606_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n290_), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n581_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n291_), .ZN(G1345gat));
  NOR2_X1   g652(.A1(new_n849_), .A2(new_n626_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT61), .B(G155gat), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  OAI21_X1  g655(.A(G162gat), .B1(new_n849_), .B2(new_n673_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n654_), .A2(G162gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n849_), .B2(new_n858_), .ZN(G1347gat));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n818_), .A2(new_n820_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n791_), .A2(new_n573_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(KEYINPUT116), .A3(new_n776_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n802_), .C1(new_n806_), .C2(new_n788_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n809_), .B1(new_n864_), .B2(new_n798_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n813_), .B1(new_n865_), .B2(new_n512_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n811_), .A2(KEYINPUT57), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n797_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n861_), .B1(new_n868_), .B2(new_n626_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n712_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n611_), .A2(new_n385_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n262_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n606_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n860_), .B1(new_n874_), .B2(new_n209_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n347_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT62), .B(G169gat), .C1(new_n873_), .C2(new_n606_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(G1348gat));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n869_), .B2(new_n712_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n647_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n581_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n872_), .A2(G176gat), .A3(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n870_), .A2(new_n883_), .A3(new_n872_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n882_), .A2(new_n884_), .B1(new_n885_), .B2(new_n207_), .ZN(G1349gat));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n871_), .A2(new_n626_), .A3(new_n262_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n880_), .A2(new_n881_), .A3(new_n888_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n889_), .A2(new_n217_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n626_), .A2(new_n229_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n826_), .A2(new_n647_), .A3(new_n872_), .A4(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n893_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n887_), .B1(new_n890_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n889_), .A2(new_n217_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n898_), .A2(KEYINPUT123), .A3(new_n895_), .A4(new_n894_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n873_), .B2(new_n673_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n512_), .A2(new_n232_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n873_), .B2(new_n902_), .ZN(G1351gat));
  AOI211_X1 g702(.A(new_n337_), .B(new_n871_), .C1(new_n815_), .C2(new_n821_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n607_), .ZN(new_n905_));
  INV_X1    g704(.A(G197gat), .ZN(new_n906_));
  OR3_X1    g705(.A1(new_n905_), .A2(KEYINPUT124), .A3(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n905_), .B2(new_n906_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n906_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n904_), .A2(new_n883_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT125), .B(G204gat), .Z(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1353gat));
  AND2_X1   g712(.A1(new_n904_), .A2(new_n547_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT63), .B(G211gat), .Z(new_n916_));
  AND3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n914_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(G1354gat));
  NAND2_X1  g719(.A1(new_n904_), .A2(new_n623_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n654_), .A2(G218gat), .ZN(new_n922_));
  AOI22_X1  g721(.A1(new_n921_), .A2(G218gat), .B1(new_n904_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1355gat));
endmodule


