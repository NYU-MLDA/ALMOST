//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT9), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G85gat), .A3(G92gat), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n204_), .A2(new_n206_), .A3(new_n211_), .A4(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n209_), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT65), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n208_), .A2(new_n210_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(KEYINPUT64), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n221_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n223_), .A2(new_n221_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n218_), .A2(new_n220_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n215_), .B1(new_n228_), .B2(new_n205_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n205_), .A2(new_n215_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT64), .B(KEYINPUT7), .ZN(new_n231_));
  MUX2_X1   g030(.A(new_n223_), .B(new_n231_), .S(new_n221_), .Z(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n232_), .B2(new_n211_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n214_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT15), .ZN(new_n235_));
  INV_X1    g034(.A(G50gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G43gat), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G50gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G36gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G29gat), .ZN(new_n244_));
  INV_X1    g043(.A(G29gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G36gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n242_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n242_), .B2(new_n249_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n235_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n249_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n250_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n242_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT15), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n234_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT35), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n264_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n251_), .A2(new_n252_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n268_), .B(new_n214_), .C1(new_n229_), .C2(new_n233_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n260_), .A2(new_n266_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n269_), .A2(new_n267_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(KEYINPUT71), .A3(new_n266_), .A4(new_n260_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n260_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n234_), .A2(new_n259_), .A3(KEYINPUT70), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n265_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G190gat), .B(G218gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G134gat), .B(G162gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT36), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n275_), .A2(new_n280_), .A3(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(KEYINPUT36), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT37), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(KEYINPUT73), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n272_), .A2(new_n274_), .B1(new_n279_), .B2(new_n265_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(new_n286_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT37), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n284_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(KEYINPUT72), .B(KEYINPUT37), .C1(new_n285_), .C2(new_n287_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n290_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT74), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n290_), .A2(new_n301_), .A3(new_n297_), .A4(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT75), .ZN(new_n305_));
  INV_X1    g104(.A(G15gat), .ZN(new_n306_));
  INV_X1    g105(.A(G22gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G15gat), .A2(G22gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G1gat), .A2(G8gat), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n308_), .A2(new_n309_), .B1(KEYINPUT14), .B2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n305_), .B(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(G57gat), .B(G64gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT11), .ZN(new_n314_));
  XOR2_X1   g113(.A(G71gat), .B(G78gat), .Z(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n314_), .A2(new_n315_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n313_), .A2(KEYINPUT11), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n312_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT76), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n320_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G127gat), .B(G155gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT16), .ZN(new_n327_));
  XOR2_X1   g126(.A(G183gat), .B(G211gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT17), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n325_), .B(new_n331_), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n330_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n323_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n303_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n234_), .A2(new_n319_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT67), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n234_), .A2(new_n319_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n319_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n341_), .B1(new_n342_), .B2(new_n337_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G120gat), .B(G148gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT5), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G176gat), .B(G204gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n353_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n345_), .A2(new_n348_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT13), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(KEYINPUT13), .A3(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n336_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT78), .ZN(new_n363_));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT83), .B1(G183gat), .B2(G190gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(G176gat), .B1(KEYINPUT84), .B2(KEYINPUT22), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G169gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n379_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(G183gat), .B2(G190gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(KEYINPUT24), .ZN(new_n391_));
  OR2_X1    g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n389_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  INV_X1    g194(.A(G190gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT26), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(G190gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(KEYINPUT82), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT26), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n396_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n384_), .B1(new_n394_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n408_));
  AND2_X1   g207(.A1(G197gat), .A2(G204gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G197gat), .A2(G204gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G211gat), .B(G218gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT21), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n412_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n409_), .A2(new_n410_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(new_n412_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n416_), .B2(KEYINPUT21), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT20), .B1(new_n407_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT22), .B(G169gat), .ZN(new_n419_));
  INV_X1    g218(.A(G176gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n390_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n378_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n386_), .B1(new_n426_), .B2(new_n379_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT91), .B1(new_n427_), .B2(new_n376_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n388_), .A2(new_n429_), .A3(new_n377_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n422_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n375_), .A2(new_n380_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n393_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n395_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT26), .B(G190gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT90), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n399_), .A2(G190gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n396_), .A2(KEYINPUT26), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT90), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n434_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n433_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n417_), .B1(new_n431_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n418_), .B1(new_n443_), .B2(KEYINPUT92), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n411_), .A2(new_n412_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n415_), .A2(new_n412_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT21), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n413_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n422_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n429_), .B1(new_n388_), .B2(new_n377_), .ZN(new_n451_));
  AOI211_X1 g250(.A(KEYINPUT91), .B(new_n376_), .C1(new_n385_), .C2(new_n387_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n437_), .A2(new_n440_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n432_), .B(new_n393_), .C1(new_n454_), .C2(new_n434_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n449_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n372_), .B1(new_n444_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n449_), .A3(new_n455_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n407_), .B2(new_n417_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n462_), .A3(new_n372_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n369_), .B1(new_n459_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n372_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n388_), .A2(new_n393_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n401_), .A2(new_n405_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n467_), .A2(new_n468_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n461_), .B1(new_n469_), .B2(new_n449_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n443_), .A2(KEYINPUT92), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n466_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n368_), .A3(new_n463_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n465_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT27), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(G155gat), .A2(G162gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G155gat), .A2(G162gat), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT2), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(KEYINPUT87), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT3), .ZN(new_n484_));
  INV_X1    g283(.A(G141gat), .ZN(new_n485_));
  INV_X1    g284(.A(G148gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n482_), .B1(new_n481_), .B2(KEYINPUT87), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n480_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT1), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n478_), .A2(new_n492_), .A3(new_n479_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n485_), .A2(new_n486_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n493_), .A2(new_n481_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(KEYINPUT29), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT28), .Z(new_n499_));
  AOI21_X1  g298(.A(new_n449_), .B1(KEYINPUT29), .B2(new_n497_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G228gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(G78gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(new_n203_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G22gat), .B(G50gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n501_), .A2(new_n502_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n444_), .A2(new_n372_), .A3(new_n458_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n460_), .A2(new_n462_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n466_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n476_), .B1(new_n515_), .B2(new_n369_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n443_), .A2(KEYINPUT92), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n458_), .A3(new_n470_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n464_), .B1(new_n518_), .B2(new_n466_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT97), .B1(new_n519_), .B2(new_n368_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n521_));
  NOR4_X1   g320(.A1(new_n459_), .A2(new_n521_), .A3(new_n369_), .A4(new_n464_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT98), .B(new_n516_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n474_), .A2(new_n521_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n473_), .A2(KEYINPUT97), .A3(new_n368_), .A4(new_n463_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT98), .B1(new_n527_), .B2(new_n516_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n477_), .B(new_n511_), .C1(new_n524_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n477_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n516_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT98), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n532_), .B1(new_n535_), .B2(new_n523_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(KEYINPUT99), .A3(new_n511_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G71gat), .B(G99gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n238_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT30), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT31), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT85), .B(G15gat), .Z(new_n543_));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n407_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n542_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT86), .ZN(new_n548_));
  XOR2_X1   g347(.A(G127gat), .B(G134gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G113gat), .B(G120gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G1gat), .B(G29gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G57gat), .B(G85gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n497_), .A2(new_n551_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G113gat), .B(G120gat), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n549_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G127gat), .B(G134gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n550_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(KEYINPUT4), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT4), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n558_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n497_), .A2(new_n551_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n558_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n557_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n570_), .A2(new_n574_), .A3(new_n557_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n548_), .A2(new_n551_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n552_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n473_), .A2(new_n463_), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n583_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT33), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n557_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n566_), .A2(new_n569_), .A3(new_n558_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n575_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n586_), .B(new_n557_), .C1(new_n570_), .C2(new_n574_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n475_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n465_), .A2(KEYINPUT94), .A3(new_n474_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n585_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n511_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT96), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n459_), .A2(new_n369_), .A3(new_n464_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n368_), .B1(new_n473_), .B2(new_n463_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n593_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n592_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n595_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n585_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n511_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n578_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n477_), .B(new_n609_), .C1(new_n524_), .C2(new_n528_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n598_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n552_), .A2(new_n579_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n538_), .A2(new_n581_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n312_), .B(new_n268_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT79), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(G229gat), .A3(G233gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n259_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(new_n312_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n312_), .A2(new_n268_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G113gat), .B(G141gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT80), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G169gat), .B(G197gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n616_), .A2(new_n621_), .A3(new_n626_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n613_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT78), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n336_), .B2(new_n361_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n363_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT100), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n363_), .A2(new_n632_), .A3(new_n637_), .A4(new_n634_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n578_), .A2(G1gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n361_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n630_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT101), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n291_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n613_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n648_), .A3(new_n335_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n578_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n640_), .A2(new_n641_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n642_), .A2(new_n650_), .A3(new_n651_), .ZN(G1324gat));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n536_), .A2(G8gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n636_), .A2(new_n638_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT102), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  OAI21_X1  g457(.A(G8gat), .B1(new_n649_), .B2(new_n536_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT39), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n658_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n654_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n663_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n653_), .A3(new_n661_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n649_), .B2(new_n612_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT41), .Z(new_n669_));
  INV_X1    g468(.A(new_n635_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n612_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n306_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(G1326gat));
  OAI21_X1  g472(.A(G22gat), .B1(new_n649_), .B2(new_n511_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT42), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(new_n307_), .A3(new_n597_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(new_n335_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n632_), .A2(new_n643_), .A3(new_n678_), .A4(new_n647_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n578_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n613_), .A2(KEYINPUT43), .A3(new_n303_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n538_), .A2(new_n581_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n611_), .A2(new_n612_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n303_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n300_), .A2(KEYINPUT105), .A3(new_n302_), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n684_), .A2(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n683_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n611_), .A2(new_n612_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n580_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n300_), .A2(KEYINPUT105), .A3(new_n302_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT105), .B1(new_n300_), .B2(new_n302_), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n692_), .A2(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n682_), .B1(new_n691_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n645_), .A2(new_n678_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT107), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n682_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n684_), .A2(new_n685_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n687_), .A2(new_n688_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n683_), .B(new_n690_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT106), .B1(new_n696_), .B2(KEYINPUT43), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707_));
  INV_X1    g506(.A(new_n699_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n700_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n691_), .A2(new_n697_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n699_), .B1(new_n712_), .B2(new_n701_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT44), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n578_), .A2(new_n245_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n681_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  NAND2_X1  g516(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n536_), .B1(new_n713_), .B2(KEYINPUT44), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n243_), .B1(new_n711_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n536_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n679_), .A2(new_n243_), .A3(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n718_), .B1(new_n720_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT110), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n718_), .B(new_n727_), .C1(new_n720_), .C2(new_n724_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n711_), .A2(new_n671_), .A3(new_n714_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G43gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n679_), .A2(new_n238_), .A3(new_n671_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(KEYINPUT47), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1330gat));
  NAND3_X1  g538(.A1(new_n679_), .A2(new_n236_), .A3(new_n597_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT111), .B1(new_n715_), .B2(new_n597_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n711_), .A2(KEYINPUT111), .A3(new_n597_), .A4(new_n714_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G50gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n741_), .B2(new_n743_), .ZN(G1331gat));
  NOR2_X1   g543(.A1(new_n613_), .A2(new_n630_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n336_), .A2(new_n643_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n578_), .B1(new_n747_), .B2(KEYINPUT112), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(KEYINPUT112), .B2(new_n747_), .ZN(new_n749_));
  INV_X1    g548(.A(G57gat), .ZN(new_n750_));
  AND4_X1   g549(.A1(new_n631_), .A2(new_n648_), .A3(new_n361_), .A4(new_n335_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n578_), .A2(new_n750_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n749_), .A2(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(G1332gat));
  INV_X1    g552(.A(G64gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n751_), .B2(new_n721_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT48), .Z(new_n756_));
  INV_X1    g555(.A(new_n747_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n754_), .A3(new_n721_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1333gat));
  NAND2_X1  g558(.A1(new_n751_), .A2(new_n671_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G71gat), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n612_), .A2(G71gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n747_), .B2(new_n763_), .ZN(G1334gat));
  AOI21_X1  g563(.A(new_n504_), .B1(new_n751_), .B2(new_n597_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT50), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n757_), .A2(new_n504_), .A3(new_n597_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1335gat));
  NAND4_X1  g567(.A1(new_n745_), .A2(new_n361_), .A3(new_n678_), .A4(new_n647_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT113), .ZN(new_n770_));
  AOI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n680_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n643_), .A2(new_n630_), .A3(new_n335_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n698_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n680_), .A2(G85gat), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT114), .Z(new_n776_));
  AOI21_X1  g575(.A(new_n771_), .B1(new_n774_), .B2(new_n776_), .ZN(G1336gat));
  INV_X1    g576(.A(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G92gat), .B1(new_n778_), .B2(new_n536_), .ZN(new_n779_));
  INV_X1    g578(.A(G92gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n770_), .A2(new_n780_), .A3(new_n721_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT115), .Z(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n778_), .B2(new_n612_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n770_), .A2(new_n671_), .A3(new_n202_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n770_), .A2(new_n203_), .A3(new_n597_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n774_), .A2(new_n597_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G106gat), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT52), .B(new_n203_), .C1(new_n774_), .C2(new_n597_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n795_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1339gat));
  NAND2_X1  g597(.A1(new_n615_), .A2(new_n619_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n619_), .B1(new_n312_), .B2(new_n268_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n626_), .B1(new_n618_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n629_), .A2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(new_n356_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n339_), .A2(KEYINPUT67), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n339_), .A2(KEYINPUT67), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n344_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n341_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(KEYINPUT55), .A3(new_n345_), .ZN(new_n810_));
  OR3_X1    g609(.A1(new_n807_), .A2(KEYINPUT55), .A3(new_n808_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n353_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT56), .B(new_n353_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n804_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n303_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT58), .B(new_n804_), .C1(new_n817_), .C2(new_n819_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n630_), .A2(new_n356_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n815_), .A2(new_n816_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n818_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n803_), .A2(new_n357_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n646_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT57), .B(new_n646_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n825_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n678_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n362_), .A2(new_n631_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT54), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n362_), .A2(new_n838_), .A3(new_n631_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n538_), .A2(new_n680_), .A3(new_n671_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(KEYINPUT118), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n834_), .A2(new_n678_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n842_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n630_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(KEYINPUT119), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(KEYINPUT119), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n841_), .A2(new_n853_), .A3(new_n843_), .A4(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT119), .B(new_n851_), .C1(new_n846_), .C2(new_n842_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n631_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n850_), .B1(new_n849_), .B2(new_n857_), .ZN(G1340gat));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n643_), .B2(G120gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n844_), .A2(new_n847_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n643_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI211_X1 g663(.A(KEYINPUT120), .B(new_n643_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G120gat), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n848_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1341gat));
  NAND3_X1  g667(.A1(new_n844_), .A2(new_n847_), .A3(new_n335_), .ZN(new_n869_));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n855_), .A2(new_n856_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n335_), .A2(G127gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT121), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n871_), .A2(new_n875_), .A3(KEYINPUT122), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1342gat));
  AOI21_X1  g679(.A(G134gat), .B1(new_n848_), .B2(new_n647_), .ZN(new_n881_));
  INV_X1    g680(.A(G134gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT123), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n882_), .A2(KEYINPUT123), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n303_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n881_), .B1(new_n872_), .B2(new_n885_), .ZN(G1343gat));
  NOR3_X1   g685(.A1(new_n846_), .A2(new_n511_), .A3(new_n671_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n721_), .A2(new_n578_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n631_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n485_), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n643_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n486_), .ZN(G1345gat));
  NOR2_X1   g692(.A1(new_n889_), .A2(new_n678_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT61), .B(G155gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(new_n889_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G162gat), .B1(new_n897_), .B2(new_n647_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n703_), .A2(G162gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(new_n899_), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n580_), .A2(new_n536_), .A3(new_n597_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n841_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G169gat), .B1(new_n902_), .B2(new_n631_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n903_), .A2(KEYINPUT62), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n630_), .A2(new_n419_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT124), .Z(new_n907_));
  OAI22_X1  g706(.A1(new_n904_), .A2(new_n905_), .B1(new_n902_), .B2(new_n907_), .ZN(G1348gat));
  NOR2_X1   g707(.A1(new_n902_), .A2(new_n643_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n420_), .ZN(G1349gat));
  NOR2_X1   g709(.A1(new_n902_), .A2(new_n678_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(G183gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n434_), .B2(new_n911_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n902_), .B2(new_n303_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n646_), .A2(new_n454_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT125), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n902_), .B2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n887_), .A2(new_n721_), .A3(new_n578_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n631_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n643_), .ZN(new_n921_));
  INV_X1    g720(.A(G204gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(KEYINPUT126), .B2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT126), .B(G204gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n921_), .B2(new_n924_), .ZN(G1353gat));
  AOI21_X1  g724(.A(new_n678_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT127), .Z(new_n927_));
  NOR2_X1   g726(.A1(new_n918_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n918_), .B2(new_n303_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n646_), .A2(G218gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n918_), .B2(new_n932_), .ZN(G1355gat));
endmodule


