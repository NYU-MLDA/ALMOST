//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G1gat), .B(G29gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT0), .ZN(new_n204_));
  INV_X1    g003(.A(G57gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT98), .B(G85gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(G141gat), .ZN(new_n212_));
  INV_X1    g011(.A(G148gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT3), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n211_), .A2(new_n214_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G155gat), .ZN(new_n220_));
  INV_X1    g019(.A(G162gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n209_), .B1(new_n219_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT84), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n229_), .A2(new_n230_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n214_), .A2(new_n211_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n216_), .A2(new_n218_), .ZN(new_n233_));
  OAI211_X1 g032(.A(KEYINPUT86), .B(new_n231_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT1), .B1(new_n223_), .B2(new_n224_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n229_), .A2(new_n237_), .A3(new_n230_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n238_), .A3(new_n222_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT85), .ZN(new_n240_));
  XOR2_X1   g039(.A(G141gat), .B(G148gat), .Z(new_n241_));
  AND3_X1   g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n235_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(new_n245_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G225gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n244_), .A2(KEYINPUT97), .A3(new_n248_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n249_), .B1(new_n244_), .B2(KEYINPUT97), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n239_), .A2(new_n241_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT85), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n257_), .A2(new_n258_), .B1(new_n226_), .B2(new_n234_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT97), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n254_), .B1(new_n255_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n253_), .B1(new_n262_), .B2(KEYINPUT4), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n244_), .A2(KEYINPUT97), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n249_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n252_), .B1(new_n266_), .B2(new_n254_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n208_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n251_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n208_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n245_), .B1(new_n266_), .B2(new_n254_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n269_), .B(new_n270_), .C1(new_n271_), .C2(new_n253_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT25), .B(G183gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G190gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT23), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n278_), .A2(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT24), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT93), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n288_), .A3(KEYINPUT24), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n282_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n291_));
  OR3_X1    g090(.A1(new_n284_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n284_), .B2(new_n290_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n285_), .B(KEYINPUT95), .Z(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT22), .B(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT96), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT96), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n296_), .A2(new_n297_), .A3(new_n303_), .A4(new_n300_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n292_), .A2(new_n293_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G197gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(G204gat), .ZN(new_n307_));
  INV_X1    g106(.A(G204gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(G197gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT21), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G218gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G211gat), .ZN(new_n312_));
  INV_X1    g111(.A(G211gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G218gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n306_), .B2(G204gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n308_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n317_), .B(new_n318_), .C1(G197gat), .C2(new_n308_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n310_), .B(new_n315_), .C1(new_n319_), .C2(KEYINPUT21), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n312_), .A2(new_n314_), .A3(KEYINPUT89), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT89), .B1(new_n312_), .B2(new_n314_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n319_), .B(KEYINPUT21), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n305_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G169gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT22), .B1(new_n326_), .B2(KEYINPUT79), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(G169gat), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n327_), .A2(new_n330_), .A3(new_n299_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n285_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n331_), .A2(new_n295_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n286_), .B2(new_n282_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n326_), .A2(new_n299_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(KEYINPUT77), .A3(KEYINPUT24), .A4(new_n285_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339_));
  NAND2_X1  g138(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT26), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT26), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT75), .A3(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G183gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT25), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G183gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n339_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n274_), .A2(KEYINPUT76), .A3(new_n341_), .A4(new_n343_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n338_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n278_), .A2(new_n280_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n282_), .A2(new_n281_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n283_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n333_), .B1(new_n352_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n324_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n325_), .A2(KEYINPUT20), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n305_), .B2(new_n324_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n361_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT18), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT32), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT99), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n324_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n320_), .A2(new_n323_), .A3(KEYINPUT91), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n284_), .A2(new_n290_), .ZN(new_n381_));
  AND4_X1   g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .A4(new_n301_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n365_), .B1(new_n382_), .B2(new_n369_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n325_), .A2(KEYINPUT20), .A3(new_n367_), .A4(new_n362_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n376_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n371_), .A2(new_n377_), .B1(KEYINPUT100), .B2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n273_), .B(new_n386_), .C1(KEYINPUT100), .C2(new_n385_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n272_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n263_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n390_), .A2(KEYINPUT33), .A3(new_n269_), .A4(new_n270_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n366_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n375_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n270_), .B1(new_n262_), .B2(new_n252_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n250_), .A2(new_n251_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n271_), .B2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n389_), .A2(new_n391_), .A3(new_n394_), .A4(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n387_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400_));
  XOR2_X1   g199(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G15gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT81), .ZN(new_n404_));
  INV_X1    g203(.A(G15gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n402_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G43gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n410_), .B(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n352_), .A2(new_n359_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n333_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n418_), .B(new_n333_), .C1(new_n352_), .C2(new_n359_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n417_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n350_), .A2(new_n351_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n338_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n283_), .B(KEYINPUT78), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n421_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n418_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n360_), .A2(new_n419_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n416_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n424_), .A2(new_n432_), .A3(new_n249_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n249_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n401_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n422_), .A2(new_n423_), .A3(new_n417_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n416_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n248_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n424_), .A2(new_n432_), .A3(new_n249_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n401_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n400_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n441_), .A3(new_n400_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n244_), .A2(KEYINPUT29), .B1(new_n379_), .B2(new_n380_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G228gat), .A2(G233gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n324_), .A2(new_n446_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n244_), .B2(KEYINPUT29), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n450_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n447_), .A2(new_n451_), .A3(new_n452_), .A4(new_n454_), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n445_), .A2(new_n446_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n449_), .A2(new_n450_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n453_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  XOR2_X1   g261(.A(G22gat), .B(G50gat), .Z(new_n463_));
  NAND3_X1  g262(.A1(new_n259_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n244_), .B2(KEYINPUT29), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  NAND3_X1  g268(.A1(new_n459_), .A2(new_n461_), .A3(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n467_), .B(new_n468_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n455_), .B(new_n458_), .C1(new_n471_), .C2(new_n460_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n443_), .A2(new_n444_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n399_), .A2(new_n473_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n470_), .A2(new_n472_), .B1(new_n441_), .B2(new_n435_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n472_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n443_), .A2(new_n444_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT27), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n375_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n481_));
  OR3_X1    g280(.A1(new_n392_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n273_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n474_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n489_));
  AND3_X1   g288(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT10), .B(G99gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(G106gat), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT9), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT64), .B(G92gat), .Z(new_n496_));
  INV_X1    g295(.A(G85gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499_));
  INV_X1    g298(.A(G92gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n501_), .B2(KEYINPUT9), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n494_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n504_), .B(new_n505_), .C1(G99gat), .C2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(G99gat), .ZN(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n507_), .B(new_n508_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(KEYINPUT67), .A3(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n510_), .A2(new_n512_), .A3(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n501_), .A2(new_n499_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT8), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n492_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n510_), .A2(KEYINPUT66), .A3(new_n492_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n501_), .A2(KEYINPUT8), .A3(new_n499_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n503_), .B1(new_n521_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n530_));
  XOR2_X1   g329(.A(G71gat), .B(G78gat), .Z(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n489_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n526_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n539_), .A2(new_n525_), .B1(new_n520_), .B2(KEYINPUT8), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT12), .B(new_n535_), .C1(new_n540_), .C2(new_n503_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n528_), .A2(new_n536_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n537_), .A2(new_n541_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n542_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n528_), .A2(new_n536_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n540_), .A2(new_n503_), .A3(new_n535_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G120gat), .B(G148gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT5), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n555_), .A2(KEYINPUT13), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n544_), .A2(new_n548_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n552_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n560_), .B2(new_n554_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n488_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G43gat), .B(G50gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G29gat), .B(G36gat), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT70), .ZN(new_n565_));
  INV_X1    g364(.A(G36gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(G29gat), .ZN(new_n567_));
  INV_X1    g366(.A(G29gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(G36gat), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n567_), .A2(new_n569_), .A3(KEYINPUT70), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n564_), .A2(KEYINPUT70), .ZN(new_n575_));
  INV_X1    g374(.A(new_n563_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G15gat), .B(G22gat), .ZN(new_n579_));
  INV_X1    g378(.A(G8gat), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G1gat), .B(G8gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n578_), .B(new_n584_), .Z(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT15), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n571_), .A2(new_n588_), .A3(new_n577_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n584_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n578_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(new_n584_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n586_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G169gat), .B(G197gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(KEYINPUT74), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT74), .B1(new_n595_), .B2(new_n599_), .ZN(new_n602_));
  OAI22_X1  g401(.A1(new_n601_), .A2(new_n602_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT13), .B1(new_n555_), .B2(new_n556_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n560_), .A2(new_n558_), .A3(new_n554_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(KEYINPUT68), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n562_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n562_), .A2(new_n603_), .A3(KEYINPUT102), .A4(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n521_), .A2(new_n527_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n503_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n578_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n589_), .A2(new_n590_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n614_), .B(new_n619_), .C1(new_n528_), .C2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n614_), .A2(KEYINPUT71), .A3(new_n619_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n617_), .A2(new_n618_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n620_), .A2(new_n528_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n528_), .A2(new_n578_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n623_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n625_), .B(new_n626_), .C1(KEYINPUT71), .C2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(KEYINPUT36), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n624_), .A2(new_n628_), .A3(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n631_), .B(KEYINPUT36), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n624_), .B2(new_n628_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT103), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n584_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(new_n536_), .ZN(new_n641_));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT16), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT17), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n641_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n647_), .B2(new_n641_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT73), .Z(new_n651_));
  NOR2_X1   g450(.A1(new_n638_), .A2(new_n651_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n487_), .A2(new_n611_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n202_), .B1(new_n653_), .B2(new_n273_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n636_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT72), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n624_), .A2(new_n628_), .A3(new_n632_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT37), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n637_), .A2(new_n656_), .A3(KEYINPUT37), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n651_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n607_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n487_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n273_), .A2(new_n202_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n654_), .B1(new_n671_), .B2(KEYINPUT38), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT104), .B(KEYINPUT38), .C1(new_n668_), .C2(new_n669_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n670_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n672_), .B(KEYINPUT105), .C1(new_n676_), .C2(new_n673_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n482_), .A2(new_n483_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n487_), .A2(new_n611_), .A3(new_n682_), .A4(new_n652_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G8gat), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT39), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT107), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n686_), .A2(new_n691_), .A3(new_n687_), .A4(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n686_), .A2(new_n688_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT39), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n690_), .A2(new_n692_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n665_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n580_), .A3(new_n682_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n695_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1325gat));
  INV_X1    g500(.A(new_n478_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n653_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G15gat), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT41), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(KEYINPUT41), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n696_), .A2(new_n405_), .A3(new_n702_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n476_), .A2(G22gat), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT110), .Z(new_n710_));
  NOR2_X1   g509(.A1(new_n665_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n653_), .A2(new_n477_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G22gat), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n715_), .B1(new_n713_), .B2(new_n714_), .ZN(G1327gat));
  NAND2_X1  g515(.A1(new_n435_), .A2(new_n441_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n476_), .A2(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n435_), .A2(new_n400_), .A3(new_n441_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n472_), .B(new_n470_), .C1(new_n719_), .C2(new_n442_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n682_), .A2(new_n273_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n721_), .A2(new_n722_), .B1(new_n399_), .B2(new_n473_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n607_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n651_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n637_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G29gat), .B1(new_n729_), .B2(new_n273_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT37), .B1(new_n637_), .B2(new_n656_), .ZN(new_n731_));
  NOR4_X1   g530(.A1(new_n633_), .A2(new_n636_), .A3(KEYINPUT72), .A4(new_n659_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT111), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n660_), .A2(new_n734_), .A3(new_n661_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n721_), .A2(new_n722_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n474_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT112), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n741_), .B(KEYINPUT43), .C1(new_n723_), .C2(new_n736_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n662_), .A2(new_n739_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n723_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n742_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n611_), .A2(new_n651_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(KEYINPUT44), .A3(new_n748_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n749_), .A2(G29gat), .A3(new_n273_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n748_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n730_), .B1(new_n750_), .B2(new_n753_), .ZN(G1328gat));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n723_), .B2(new_n736_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n744_), .B1(new_n755_), .B2(KEYINPUT112), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n747_), .B1(new_n756_), .B2(new_n742_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n484_), .B1(new_n757_), .B2(KEYINPUT44), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n566_), .B1(new_n758_), .B2(new_n753_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n728_), .A2(G36gat), .A3(new_n484_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT45), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT113), .B(KEYINPUT46), .Z(new_n762_));
  NOR3_X1   g561(.A1(new_n759_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n762_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n749_), .A2(new_n682_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT44), .B1(new_n746_), .B2(new_n748_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G36gat), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n761_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n763_), .A2(new_n769_), .ZN(G1329gat));
  OAI21_X1  g569(.A(new_n413_), .B1(new_n728_), .B2(new_n478_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT114), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n749_), .A2(G43gat), .A3(new_n717_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n766_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g574(.A(G50gat), .B1(new_n729_), .B2(new_n477_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n749_), .A2(G50gat), .A3(new_n477_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n753_), .ZN(G1331gat));
  NAND2_X1  g577(.A1(new_n562_), .A2(new_n606_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n595_), .A2(new_n599_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n602_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n600_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n723_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n652_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G57gat), .B1(new_n785_), .B2(new_n485_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n779_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n787_), .A2(new_n662_), .A3(new_n651_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n788_), .A2(KEYINPUT115), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(KEYINPUT115), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n782_), .A3(new_n487_), .A4(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT116), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n273_), .A2(new_n205_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n786_), .B1(new_n792_), .B2(new_n793_), .ZN(G1332gat));
  OAI21_X1  g593(.A(G64gat), .B1(new_n785_), .B2(new_n484_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT48), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n484_), .A2(G64gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n792_), .B2(new_n797_), .ZN(G1333gat));
  OR2_X1    g597(.A1(new_n478_), .A2(G71gat), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n784_), .A2(new_n702_), .A3(new_n652_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G71gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n800_), .A3(G71gat), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI22_X1  g603(.A1(new_n792_), .A2(new_n799_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT117), .ZN(G1334gat));
  OAI21_X1  g605(.A(G78gat), .B1(new_n785_), .B2(new_n476_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT50), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n476_), .A2(G78gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n792_), .B2(new_n809_), .ZN(G1335gat));
  NAND2_X1  g609(.A1(new_n784_), .A2(new_n727_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n497_), .A3(new_n273_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n783_), .A2(new_n725_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n746_), .A2(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n815_), .A2(KEYINPUT118), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(KEYINPUT118), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n485_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n813_), .B1(new_n818_), .B2(new_n497_), .ZN(G1336gat));
  OAI21_X1  g618(.A(new_n500_), .B1(new_n811_), .B2(new_n484_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT119), .Z(new_n821_));
  NOR2_X1   g620(.A1(new_n816_), .A2(new_n817_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n484_), .A2(new_n496_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n822_), .B2(new_n823_), .ZN(G1337gat));
  NOR2_X1   g623(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n493_), .B(new_n811_), .C1(new_n441_), .C2(new_n435_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n746_), .A2(new_n702_), .A3(new_n814_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(G99gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n825_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1338gat));
  NAND3_X1  g631(.A1(new_n812_), .A2(new_n508_), .A3(new_n477_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n746_), .A2(new_n477_), .A3(new_n814_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(new_n835_), .A3(G106gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n834_), .B2(G106gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n833_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT53), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n833_), .B(new_n840_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1339gat));
  NAND2_X1  g641(.A1(new_n484_), .A2(new_n273_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n718_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT122), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n599_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n593_), .B2(new_n586_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n554_), .B(new_n847_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n537_), .A2(new_n543_), .A3(new_n541_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT55), .A3(new_n542_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n544_), .A2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n850_), .B(new_n852_), .C1(new_n542_), .C2(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n552_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n848_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n858_), .A2(KEYINPUT58), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n731_), .A2(new_n732_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n858_), .B2(KEYINPUT58), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n857_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n603_), .A3(new_n554_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n847_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n555_), .A2(new_n556_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n637_), .B1(new_n864_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n862_), .B1(KEYINPUT57), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(KEYINPUT57), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n725_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n603_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n663_), .A2(new_n874_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n875_), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT121), .B1(new_n875_), .B2(KEYINPUT54), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n875_), .A2(KEYINPUT54), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n845_), .B1(new_n873_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(G113gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n603_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n873_), .B2(new_n879_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n880_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n872_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n651_), .B1(new_n870_), .B2(new_n888_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n877_), .A2(new_n878_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n876_), .B2(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n891_), .B(new_n845_), .C1(new_n884_), .C2(KEYINPUT59), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n782_), .B1(new_n887_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n883_), .B1(new_n893_), .B2(new_n882_), .ZN(G1340gat));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895_));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n779_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n881_), .A2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n787_), .B1(new_n887_), .B2(new_n892_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n896_), .ZN(G1341gat));
  INV_X1    g700(.A(G127gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n881_), .A2(new_n902_), .A3(new_n725_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n651_), .B1(new_n887_), .B2(new_n892_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n902_), .ZN(G1342gat));
  AOI21_X1  g704(.A(G134gat), .B1(new_n881_), .B2(new_n638_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n887_), .A2(new_n892_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT124), .B(G134gat), .Z(new_n908_));
  NOR2_X1   g707(.A1(new_n860_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n906_), .B1(new_n907_), .B2(new_n909_), .ZN(G1343gat));
  INV_X1    g709(.A(new_n720_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n843_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n891_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n603_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT125), .B(G141gat), .Z(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n915_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n913_), .A2(new_n603_), .A3(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n913_), .A2(new_n779_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G148gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n913_), .A2(new_n213_), .A3(new_n779_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1345gat));
  NAND4_X1  g722(.A1(new_n891_), .A2(new_n725_), .A3(new_n911_), .A4(new_n912_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1346gat));
  AOI21_X1  g725(.A(G162gat), .B1(new_n913_), .B2(new_n638_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n736_), .A2(new_n221_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n913_), .B2(new_n928_), .ZN(G1347gat));
  NOR4_X1   g728(.A1(new_n484_), .A2(new_n477_), .A3(new_n478_), .A4(new_n273_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n891_), .A2(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931_), .B2(new_n782_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  OAI211_X1 g733(.A(KEYINPUT62), .B(G169gat), .C1(new_n931_), .C2(new_n782_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n931_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n936_), .A2(new_n603_), .A3(new_n298_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n934_), .A2(new_n935_), .A3(new_n937_), .ZN(G1348gat));
  NOR2_X1   g737(.A1(new_n931_), .A2(new_n787_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(KEYINPUT126), .A3(new_n299_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT126), .B(G176gat), .Z(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n939_), .B2(new_n941_), .ZN(G1349gat));
  NOR2_X1   g741(.A1(new_n931_), .A2(new_n651_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n274_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n944_), .B1(new_n345_), .B2(new_n943_), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n931_), .B2(new_n860_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n638_), .A2(new_n275_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n931_), .B2(new_n947_), .ZN(G1351gat));
  NOR2_X1   g747(.A1(new_n484_), .A2(new_n273_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n891_), .A2(new_n603_), .A3(new_n911_), .A4(new_n949_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g750(.A(new_n787_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n891_), .A2(new_n911_), .A3(new_n949_), .A4(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n954_));
  XOR2_X1   g753(.A(new_n953_), .B(new_n954_), .Z(G1353gat));
  AOI21_X1  g754(.A(new_n651_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n891_), .A2(new_n911_), .A3(new_n949_), .A4(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  XOR2_X1   g757(.A(new_n957_), .B(new_n958_), .Z(G1354gat));
  AND2_X1   g758(.A1(new_n891_), .A2(new_n911_), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n960_), .A2(new_n311_), .A3(new_n638_), .A4(new_n949_), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n960_), .A2(new_n662_), .A3(new_n949_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n962_), .B2(new_n311_), .ZN(G1355gat));
endmodule


