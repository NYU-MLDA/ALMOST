//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n206_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n202_), .B(new_n205_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n207_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n211_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n218_), .B(new_n220_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT81), .B1(new_n223_), .B2(new_n224_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n215_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(G113gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(G113gat), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n232_), .A2(G120gat), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(G120gat), .B1(new_n232_), .B2(new_n233_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n230_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT31), .B(G43gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT83), .B(G15gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n240_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n241_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n241_), .B2(new_n245_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G57gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G85gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(G1gat), .B(G29gat), .Z(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n231_), .B(G113gat), .ZN(new_n253_));
  INV_X1    g052(.A(G120gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n232_), .A2(G120gat), .A3(new_n233_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n260_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(G141gat), .ZN(new_n262_));
  INV_X1    g061(.A(G148gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n259_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n261_), .B(new_n264_), .C1(KEYINPUT1), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(KEYINPUT84), .A3(new_n259_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n273_));
  OR3_X1    g072(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  AND4_X1   g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n267_), .B1(new_n271_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n257_), .A2(new_n258_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT90), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT90), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n267_), .B(new_n281_), .C1(new_n271_), .C2(new_n277_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n236_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n278_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(new_n257_), .A3(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT91), .B1(new_n286_), .B2(KEYINPUT4), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT91), .ZN(new_n288_));
  AOI211_X1 g087(.A(new_n288_), .B(new_n258_), .C1(new_n283_), .C2(new_n285_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n279_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G225gat), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n286_), .A2(new_n292_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n252_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n252_), .ZN(new_n297_));
  AOI211_X1 g096(.A(new_n297_), .B(new_n294_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n248_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G22gat), .B(G50gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n284_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n278_), .B2(KEYINPUT29), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n302_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n302_), .A3(new_n307_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G78gat), .B(G106gat), .Z(new_n312_));
  OR2_X1    g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G228gat), .ZN(new_n314_));
  INV_X1    g113(.A(G233gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G211gat), .B(G218gat), .Z(new_n317_));
  XOR2_X1   g116(.A(G197gat), .B(G204gat), .Z(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(KEYINPUT21), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n320_));
  INV_X1    g119(.A(G197gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(G204gat), .ZN(new_n322_));
  INV_X1    g121(.A(G204gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n322_), .A2(new_n324_), .B1(new_n321_), .B2(G204gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n325_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(KEYINPUT21), .A3(new_n317_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT87), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n316_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n333_), .B(new_n331_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n311_), .B1(KEYINPUT88), .B2(new_n312_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n313_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n313_), .B2(new_n338_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT18), .B(G64gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT19), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n205_), .A2(new_n202_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n214_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n220_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n352_));
  OAI221_X1 g151(.A(new_n332_), .B1(new_n350_), .B2(new_n351_), .C1(new_n225_), .C2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n229_), .B2(new_n331_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n349_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n325_), .A2(new_n326_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n317_), .A2(new_n357_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n358_), .B(new_n215_), .C1(new_n228_), .C2(new_n227_), .ZN(new_n359_));
  OAI22_X1  g158(.A1(new_n352_), .A2(new_n225_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n354_), .B1(new_n331_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(new_n348_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n346_), .B1(new_n356_), .B2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n355_), .B(new_n349_), .C1(new_n331_), .C2(new_n360_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT89), .B1(new_n362_), .B2(new_n348_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  AOI211_X1 g166(.A(new_n367_), .B(new_n349_), .C1(new_n359_), .C2(new_n361_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n365_), .B(new_n345_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(KEYINPUT27), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT92), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n365_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n346_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n369_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n371_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  AOI211_X1 g175(.A(KEYINPUT92), .B(KEYINPUT27), .C1(new_n373_), .C2(new_n369_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n341_), .B(new_n370_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT94), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n364_), .A2(KEYINPUT27), .A3(new_n369_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n373_), .A2(new_n369_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT92), .B1(new_n381_), .B2(KEYINPUT27), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT94), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n341_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n300_), .B1(new_n379_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT93), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n339_), .A2(new_n340_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n370_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n299_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n384_), .A2(KEYINPUT93), .A3(new_n299_), .A4(new_n389_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n291_), .B(new_n279_), .C1(new_n287_), .C2(new_n289_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n286_), .A2(new_n292_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n394_), .A2(new_n252_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT33), .B1(new_n296_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n294_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n252_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n381_), .A3(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n356_), .B2(new_n363_), .ZN(new_n403_));
  OAI221_X1 g202(.A(new_n403_), .B1(new_n372_), .B2(new_n402_), .C1(new_n296_), .C2(new_n298_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n392_), .B(new_n393_), .C1(new_n405_), .C2(new_n389_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n248_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n387_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G169gat), .B(G197gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n411_), .A2(G113gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(G113gat), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n412_), .A2(G141gat), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(G141gat), .B1(new_n412_), .B2(new_n413_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G229gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G15gat), .B(G22gat), .ZN(new_n420_));
  INV_X1    g219(.A(G1gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G8gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(G29gat), .A2(G36gat), .ZN(new_n427_));
  INV_X1    g226(.A(G43gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G29gat), .A2(G36gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(G29gat), .A2(G36gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G29gat), .A2(G36gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(G43gat), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G50gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(new_n433_), .A3(G50gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n426_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n426_), .A2(new_n438_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n419_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT15), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n430_), .A2(new_n433_), .A3(G50gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(G50gat), .B1(new_n430_), .B2(new_n433_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(KEYINPUT15), .A3(new_n437_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n426_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n440_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n418_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n417_), .A2(new_n441_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n417_), .B1(new_n441_), .B2(new_n450_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G120gat), .B(G148gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(new_n323_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT5), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(new_n204_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT71), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G230gat), .A2(G233gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT67), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  OR3_X1    g267(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n469_), .A2(new_n472_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n468_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT67), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n462_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n473_), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT10), .B(G99gat), .Z(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n487_));
  AND2_X1   g286(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT9), .ZN(new_n490_));
  AND2_X1   g289(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n487_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n486_), .B1(new_n494_), .B2(new_n466_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n468_), .B(new_n475_), .C1(new_n477_), .C2(KEYINPUT8), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n482_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(G57gat), .A2(G64gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G57gat), .A2(G64gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT11), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G57gat), .ZN(new_n501_));
  INV_X1    g300(.A(G64gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G57gat), .A2(G64gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G71gat), .ZN(new_n507_));
  INV_X1    g306(.A(G78gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G71gat), .A2(G78gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n500_), .A2(new_n506_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n513_));
  OAI221_X1 g312(.A(KEYINPUT11), .B1(new_n498_), .B2(new_n499_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n516_), .A3(new_n514_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n460_), .B1(new_n497_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT70), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT12), .B1(new_n497_), .B2(new_n520_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n497_), .A2(new_n520_), .A3(KEYINPUT12), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n460_), .C1(new_n497_), .C2(new_n520_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .A4(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n482_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n519_), .A3(new_n518_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n497_), .A2(new_n520_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(G230gat), .A3(G233gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n459_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n528_), .A2(new_n533_), .A3(new_n458_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n459_), .A2(new_n534_), .A3(KEYINPUT72), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT13), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(KEYINPUT13), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n408_), .A2(new_n454_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT75), .B1(new_n497_), .B2(new_n447_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT73), .Z(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT34), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n546_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n497_), .A2(new_n447_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT74), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n438_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n529_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n529_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT75), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(KEYINPUT35), .A3(new_n550_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT74), .B1(new_n497_), .B2(new_n447_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n497_), .A2(new_n438_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n559_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n560_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT76), .B(G134gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G162gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n551_), .A2(new_n547_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n568_), .A2(new_n575_), .A3(new_n576_), .A4(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n560_), .A2(new_n567_), .A3(new_n576_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n579_), .A2(KEYINPUT77), .A3(new_n574_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT77), .B1(new_n579_), .B2(new_n574_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT78), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n584_), .B(new_n578_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n583_), .A2(KEYINPUT37), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT37), .B1(new_n583_), .B2(new_n585_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n520_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n426_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT16), .B(G183gat), .ZN(new_n593_));
  INV_X1    g392(.A(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n592_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(new_n591_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT79), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n588_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n545_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n421_), .A3(new_n391_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT38), .ZN(new_n606_));
  INV_X1    g405(.A(new_n582_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n545_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n299_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n384_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n545_), .A2(new_n422_), .A3(new_n612_), .A4(new_n603_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT95), .Z(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n609_), .B2(new_n384_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT39), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n617_), .B(G8gat), .C1(new_n609_), .C2(new_n384_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n619_), .A3(KEYINPUT40), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1325gat));
  OAI21_X1  g423(.A(G15gat), .B1(new_n609_), .B2(new_n407_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT41), .Z(new_n626_));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n604_), .A2(new_n627_), .A3(new_n248_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n341_), .B(KEYINPUT96), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n604_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n631_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n609_), .B2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT42), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(KEYINPUT42), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT97), .B(new_n632_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1327gat));
  NAND2_X1  g440(.A1(new_n602_), .A2(new_n607_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT99), .Z(new_n643_));
  AND2_X1   g442(.A1(new_n545_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n391_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n544_), .A2(new_n601_), .A3(new_n454_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n393_), .A2(new_n392_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n389_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n407_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n387_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n647_), .B1(new_n652_), .B2(new_n588_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT37), .ZN(new_n654_));
  INV_X1    g453(.A(new_n581_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n579_), .A2(KEYINPUT77), .A3(new_n574_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n584_), .B1(new_n657_), .B2(new_n578_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n585_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n583_), .A2(KEYINPUT37), .A3(new_n585_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n408_), .A2(KEYINPUT43), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n646_), .B1(new_n653_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(KEYINPUT98), .A2(KEYINPUT44), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n665_), .A3(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n652_), .A2(new_n647_), .A3(new_n588_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n408_), .B2(new_n662_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(new_n666_), .A3(new_n667_), .A4(new_n646_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n299_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n645_), .B1(new_n674_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n545_), .A2(new_n676_), .A3(new_n612_), .A4(new_n643_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT45), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n384_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n676_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT46), .B(new_n678_), .C1(new_n679_), .C2(new_n676_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  AOI211_X1 g483(.A(new_n428_), .B(new_n407_), .C1(new_n669_), .C2(new_n673_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G43gat), .B1(new_n644_), .B2(new_n248_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT47), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n669_), .A2(new_n673_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(G43gat), .A3(new_n248_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690_));
  INV_X1    g489(.A(new_n686_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n687_), .A2(new_n692_), .ZN(G1330gat));
  AOI21_X1  g492(.A(G50gat), .B1(new_n644_), .B2(new_n631_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n435_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n389_), .ZN(G1331gat));
  INV_X1    g495(.A(new_n454_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n408_), .A2(new_n697_), .A3(new_n543_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n603_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n501_), .A3(new_n391_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n608_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n299_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT100), .ZN(G1332gat));
  OAI21_X1  g503(.A(G64gat), .B1(new_n701_), .B2(new_n384_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT48), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n699_), .A2(new_n502_), .A3(new_n612_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1333gat));
  OAI21_X1  g507(.A(G71gat), .B1(new_n701_), .B2(new_n407_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT101), .B(KEYINPUT49), .Z(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT102), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n709_), .B(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n699_), .A2(new_n507_), .A3(new_n248_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1334gat));
  NAND3_X1  g513(.A1(new_n699_), .A2(new_n508_), .A3(new_n631_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n701_), .A2(new_n633_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n716_), .A2(KEYINPUT103), .A3(new_n508_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT103), .B1(new_n716_), .B2(new_n508_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(KEYINPUT50), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT50), .B1(new_n717_), .B2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n719_), .B2(new_n720_), .ZN(G1335gat));
  AND2_X1   g520(.A1(new_n698_), .A2(new_n643_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n391_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n544_), .A2(new_n602_), .A3(new_n454_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT104), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n672_), .A2(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n299_), .A2(new_n492_), .A3(new_n491_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT105), .Z(G1336gat));
  AOI21_X1  g528(.A(G92gat), .B1(new_n722_), .B2(new_n612_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT106), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n384_), .A2(new_n489_), .A3(new_n488_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT107), .Z(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n726_), .B2(new_n733_), .ZN(G1337gat));
  AND3_X1   g533(.A1(new_n722_), .A2(new_n484_), .A3(new_n248_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n726_), .A2(new_n248_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G99gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n722_), .A2(new_n485_), .A3(new_n389_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n672_), .A2(new_n725_), .A3(new_n389_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G106gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT53), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(new_n740_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1339gat));
  INV_X1    g548(.A(G113gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n697_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n601_), .B(new_n751_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n662_), .A2(KEYINPUT54), .A3(new_n601_), .A4(new_n751_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n528_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n524_), .A2(new_n530_), .A3(new_n525_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(G230gat), .A3(G233gat), .ZN(new_n761_));
  INV_X1    g560(.A(new_n525_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(new_n523_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(KEYINPUT55), .A3(new_n522_), .A4(new_n527_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n761_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n459_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n697_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT109), .B1(new_n765_), .B2(new_n459_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n538_), .B1(new_n770_), .B2(KEYINPUT56), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n757_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n766_), .A2(new_n767_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n454_), .B1(new_n770_), .B2(KEYINPUT56), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT110), .A4(new_n538_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n448_), .A2(new_n449_), .A3(new_n419_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n418_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n416_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT111), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n416_), .A2(new_n778_), .A3(new_n779_), .A4(new_n782_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n781_), .A2(new_n451_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n540_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n772_), .A2(new_n777_), .A3(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n786_), .A2(KEYINPUT57), .A3(new_n582_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT57), .B1(new_n786_), .B2(new_n582_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n774_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n766_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n784_), .A2(new_n793_), .A3(new_n538_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n528_), .A2(new_n533_), .A3(new_n458_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n781_), .A2(new_n451_), .A3(new_n783_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT112), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n765_), .A2(new_n789_), .A3(new_n774_), .A4(new_n459_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n792_), .A2(new_n798_), .A3(KEYINPUT58), .A4(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n804_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n787_), .A2(new_n788_), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n756_), .B1(new_n806_), .B2(new_n601_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n379_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n386_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n807_), .A2(new_n391_), .A3(new_n811_), .A4(new_n248_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n750_), .B1(new_n812_), .B2(new_n454_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n754_), .A2(new_n755_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n786_), .A2(new_n582_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n588_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n786_), .A2(KEYINPUT57), .A3(new_n582_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n818_), .B1(new_n824_), .B2(new_n602_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n825_), .A2(new_n299_), .A3(new_n810_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n817_), .B1(new_n826_), .B2(new_n248_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n812_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n816_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n248_), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(KEYINPUT116), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n454_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n815_), .B1(new_n835_), .B2(G113gat), .ZN(G1340gat));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n544_), .A3(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT117), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n832_), .A2(new_n833_), .A3(new_n839_), .A4(new_n544_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(G120gat), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n812_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n254_), .B1(new_n543_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n842_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n254_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n842_), .B2(new_n601_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT118), .A2(G127gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G127gat), .B1(new_n602_), .B2(KEYINPUT118), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n846_), .B1(new_n848_), .B2(new_n849_), .ZN(G1342gat));
  AOI21_X1  g649(.A(G134gat), .B1(new_n842_), .B2(new_n607_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n662_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n825_), .A2(new_n299_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n390_), .A2(new_n248_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT119), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(new_n858_), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT120), .B(G141gat), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n860_), .A2(new_n697_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(new_n697_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1344gat));
  AOI21_X1  g663(.A(new_n543_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT121), .B(G148gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1345gat));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n860_), .A2(new_n601_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n860_), .B2(new_n601_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  AOI21_X1  g670(.A(G162gat), .B1(new_n860_), .B2(new_n607_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n662_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(G162gat), .B2(new_n873_), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n300_), .A2(new_n384_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n825_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n633_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n697_), .A3(new_n203_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n877_), .A2(KEYINPUT122), .A3(new_n697_), .A4(new_n633_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n807_), .A2(new_n697_), .A3(new_n633_), .A4(new_n875_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(new_n885_), .A3(G169gat), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n881_), .B1(new_n887_), .B2(new_n888_), .ZN(G1348gat));
  AND4_X1   g688(.A1(G176gat), .A2(new_n877_), .A3(new_n544_), .A4(new_n341_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n880_), .A2(new_n544_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n204_), .ZN(G1349gat));
  NOR3_X1   g691(.A1(new_n756_), .A2(new_n602_), .A3(new_n389_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G183gat), .B1(new_n893_), .B2(new_n875_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n878_), .B(KEYINPUT123), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n602_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n221_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n894_), .B1(new_n896_), .B2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n895_), .B2(new_n662_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n880_), .A2(new_n607_), .A3(new_n222_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1351gat));
  NAND3_X1  g700(.A1(new_n807_), .A2(new_n389_), .A3(new_n407_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(new_n391_), .A3(new_n384_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n697_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n544_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(KEYINPUT124), .B2(G204gat), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT124), .B(G204gat), .Z(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(G1353gat));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n601_), .B1(new_n910_), .B2(new_n594_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT125), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n903_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n594_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1354gat));
  AOI21_X1  g714(.A(G218gat), .B1(new_n903_), .B2(new_n607_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n588_), .A2(G218gat), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT126), .Z(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n903_), .B2(new_n918_), .ZN(G1355gat));
endmodule


