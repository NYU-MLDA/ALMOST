//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT90), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n210_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT91), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n219_), .B(new_n220_), .C1(new_n221_), .C2(new_n210_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n205_), .B(new_n206_), .C1(new_n217_), .C2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n214_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G127gat), .B(G134gat), .Z(new_n225_));
  XOR2_X1   g024(.A(G113gat), .B(G120gat), .Z(new_n226_));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n225_), .B(new_n226_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(new_n227_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n224_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n224_), .A2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT4), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n228_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n214_), .A2(new_n223_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n224_), .A2(new_n229_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n234_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT0), .ZN(new_n247_));
  INV_X1    g046(.A(G57gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G85gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n241_), .A2(new_n251_), .A3(new_n244_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n256_));
  AND2_X1   g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n257_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(G183gat), .B2(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G176gat), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT84), .B1(new_n266_), .B2(KEYINPUT22), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n265_), .B(new_n267_), .C1(new_n268_), .C2(KEYINPUT84), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n261_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n264_), .B(KEYINPUT24), .C1(G169gat), .C2(G176gat), .ZN(new_n271_));
  NOR3_X1   g070(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n257_), .A2(new_n259_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT81), .B1(new_n276_), .B2(G190gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT25), .B(G183gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G190gat), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n277_), .B(new_n278_), .C1(new_n279_), .C2(KEYINPUT81), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n271_), .A2(new_n273_), .A3(new_n275_), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n270_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G197gat), .B(G204gat), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT93), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n284_), .A2(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n290_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n282_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n264_), .B(KEYINPUT97), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n268_), .A2(new_n265_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n275_), .B1(G183gat), .B2(G190gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT96), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT96), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n302_), .B(new_n303_), .C1(G169gat), .C2(G176gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n272_), .B1(new_n279_), .B2(new_n278_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n260_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n300_), .A2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n295_), .B(new_n296_), .C1(new_n294_), .C2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT19), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT20), .B1(new_n282_), .B2(new_n294_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT95), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT98), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n300_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n297_), .A2(KEYINPUT98), .A3(new_n298_), .A4(new_n299_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n306_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n294_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n319_), .B(KEYINPUT20), .C1(new_n282_), .C2(new_n294_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n313_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n311_), .B1(new_n321_), .B2(new_n310_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G8gat), .B(G36gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT18), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G64gat), .ZN(new_n325_));
  INV_X1    g124(.A(G92gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT32), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n310_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT20), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n282_), .B2(new_n294_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(new_n317_), .B2(new_n294_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT99), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT99), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n333_), .B(new_n336_), .C1(new_n317_), .C2(new_n294_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n321_), .A2(new_n310_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n255_), .B(new_n330_), .C1(new_n340_), .C2(new_n329_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT33), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n253_), .A2(KEYINPUT100), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT100), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n251_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n345_), .B2(KEYINPUT33), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n235_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n251_), .B1(new_n243_), .B2(new_n234_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n253_), .B2(new_n342_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n327_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n340_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n338_), .A2(new_n339_), .A3(new_n327_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n341_), .B1(new_n347_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G15gat), .B(G43gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT85), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n270_), .A2(KEYINPUT30), .A3(new_n281_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT30), .B1(new_n270_), .B2(new_n281_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT86), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n360_), .B(new_n361_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n371_), .B(KEYINPUT86), .C1(new_n365_), .C2(new_n364_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT88), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n230_), .A2(KEYINPUT31), .A3(new_n228_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT31), .B1(new_n230_), .B2(new_n228_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n373_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(KEYINPUT88), .A3(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n372_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT89), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n370_), .A2(new_n372_), .A3(new_n383_), .A4(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n370_), .A2(new_n372_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n375_), .A2(new_n376_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT94), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n237_), .A2(KEYINPUT29), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n294_), .A2(KEYINPUT92), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n224_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G22gat), .B(G50gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT28), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n237_), .A2(KEYINPUT29), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n397_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n393_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n395_), .A2(new_n398_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n293_), .A2(new_n292_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(new_n291_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n397_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .A4(new_n392_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n403_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n403_), .B1(new_n402_), .B2(new_n409_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n391_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(new_n390_), .A3(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n388_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n356_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT103), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n353_), .A2(new_n354_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  AOI211_X1 g221(.A(KEYINPUT103), .B(KEYINPUT27), .C1(new_n353_), .C2(new_n354_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n354_), .A2(KEYINPUT102), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n322_), .B2(new_n352_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(KEYINPUT102), .B2(new_n354_), .ZN(new_n426_));
  OAI22_X1  g225(.A1(new_n422_), .A2(new_n423_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n413_), .A2(new_n415_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n388_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n381_), .A2(KEYINPUT89), .B1(new_n385_), .B2(new_n386_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n416_), .A2(new_n430_), .A3(new_n384_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n255_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n418_), .B1(new_n427_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT10), .B(G99gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT64), .B(G106gat), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G85gat), .B(G92gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT9), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(G85gat), .A3(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT6), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT8), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT68), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT67), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT6), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n449_), .A2(new_n451_), .A3(new_n443_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n443_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n447_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n443_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n450_), .A2(KEYINPUT6), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n448_), .A2(KEYINPUT67), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n451_), .A3(new_n443_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT68), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT65), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n454_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n439_), .B(KEYINPUT66), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n446_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n444_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n466_), .A2(new_n468_), .A3(new_n446_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n445_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G29gat), .B(G36gat), .Z(new_n471_));
  XOR2_X1   g270(.A(G43gat), .B(G50gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT15), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G232gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT34), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n473_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n475_), .B(new_n480_), .C1(new_n470_), .C2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n478_), .A2(new_n479_), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n483_), .B(KEYINPUT75), .Z(new_n484_));
  XNOR2_X1  g283(.A(new_n482_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G190gat), .B(G218gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G134gat), .B(G162gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(KEYINPUT36), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n488_), .A2(KEYINPUT36), .ZN(new_n490_));
  OR3_X1    g289(.A1(new_n485_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n489_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n435_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT104), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G57gat), .B(G64gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT69), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n496_), .A2(KEYINPUT69), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT11), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(KEYINPUT69), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G71gat), .B(G78gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n498_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n497_), .A2(KEYINPUT11), .A3(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(new_n445_), .C1(new_n467_), .C2(new_n469_), .ZN(new_n508_));
  INV_X1    g307(.A(G230gat), .ZN(new_n509_));
  INV_X1    g308(.A(G233gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n505_), .A2(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n470_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT70), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT12), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  AOI211_X1 g318(.A(KEYINPUT70), .B(new_n519_), .C1(new_n470_), .C2(new_n515_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n514_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT71), .ZN(new_n522_));
  INV_X1    g321(.A(new_n516_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n508_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n511_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n514_), .C1(new_n518_), .C2(new_n520_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n522_), .A2(new_n525_), .A3(new_n527_), .A4(new_n533_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(KEYINPUT73), .A3(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(KEYINPUT13), .A3(new_n540_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545_));
  INV_X1    g344(.A(G8gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G1gat), .B(G8gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n473_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT78), .ZN(new_n552_));
  INV_X1    g351(.A(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n474_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT79), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT79), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n559_), .A3(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n481_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n552_), .A2(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n562_), .A2(new_n556_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n558_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G169gat), .B(G197gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT80), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n558_), .A2(new_n563_), .A3(new_n560_), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n507_), .B(new_n553_), .ZN(new_n573_));
  AND2_X1   g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n574_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(KEYINPUT76), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(G183gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G211gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT77), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(KEYINPUT76), .B2(new_n578_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n578_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n583_), .B(KEYINPUT17), .Z(new_n588_));
  AOI22_X1  g387(.A1(new_n579_), .A2(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n543_), .A2(new_n544_), .A3(new_n572_), .A4(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n494_), .B1(new_n495_), .B2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n495_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n202_), .B1(new_n593_), .B2(new_n255_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT105), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n426_), .A2(new_n424_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n354_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n327_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n421_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT103), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n420_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n596_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n255_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n602_), .A2(new_n603_), .B1(new_n356_), .B2(new_n417_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n493_), .B(KEYINPUT37), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n589_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n543_), .A2(new_n544_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n572_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n202_), .A3(new_n255_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT38), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n595_), .A2(new_n615_), .ZN(G1324gat));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n546_), .A3(new_n427_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n591_), .A2(new_n592_), .A3(new_n427_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT106), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT106), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n591_), .A2(new_n592_), .A3(new_n621_), .A4(new_n427_), .ZN(new_n622_));
  AND4_X1   g421(.A1(new_n618_), .A2(new_n620_), .A3(G8gat), .A4(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n546_), .B1(new_n619_), .B2(KEYINPUT106), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n618_), .B1(new_n624_), .B2(new_n622_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n617_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT40), .B(new_n617_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  NAND2_X1  g429(.A1(new_n593_), .A2(new_n388_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G15gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  INV_X1    g432(.A(new_n388_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n612_), .A2(G15gat), .A3(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n416_), .B(KEYINPUT107), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n593_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT42), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n613_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1327gat));
  NOR2_X1   g442(.A1(new_n589_), .A2(new_n493_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT110), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n611_), .A2(new_n435_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT111), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT111), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n611_), .A2(new_n648_), .A3(new_n435_), .A4(new_n645_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n255_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT43), .B1(new_n604_), .B2(new_n605_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n435_), .A2(new_n653_), .A3(new_n606_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n609_), .A2(new_n610_), .A3(new_n589_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(KEYINPUT44), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n655_), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n656_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(G29gat), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n433_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT44), .B1(new_n655_), .B2(new_n656_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n651_), .B1(new_n664_), .B2(new_n667_), .ZN(G1328gat));
  OAI21_X1  g467(.A(new_n427_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n665_), .B(KEYINPUT108), .ZN(new_n670_));
  OAI21_X1  g469(.A(G36gat), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G36gat), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n647_), .A2(new_n672_), .A3(new_n427_), .A4(new_n649_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT45), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(KEYINPUT46), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n657_), .A2(new_n658_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n602_), .B1(new_n677_), .B2(new_n660_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n672_), .B1(new_n667_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n673_), .B(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n676_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n675_), .A2(new_n682_), .ZN(G1329gat));
  NAND2_X1  g482(.A1(new_n650_), .A2(new_n388_), .ZN(new_n684_));
  INV_X1    g483(.A(G43gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(G43gat), .B(new_n388_), .C1(new_n659_), .C2(new_n661_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(new_n670_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT47), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n686_), .B(new_n690_), .C1(new_n687_), .C2(new_n670_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1330gat));
  AOI21_X1  g491(.A(G50gat), .B1(new_n650_), .B2(new_n639_), .ZN(new_n693_));
  INV_X1    g492(.A(G50gat), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n662_), .A2(new_n694_), .A3(new_n428_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(new_n667_), .ZN(G1331gat));
  NOR2_X1   g495(.A1(new_n607_), .A2(new_n572_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n435_), .A2(new_n493_), .A3(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(KEYINPUT113), .A3(new_n609_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT113), .B1(new_n698_), .B2(new_n609_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n700_), .A2(new_n433_), .A3(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n609_), .A2(new_n589_), .A3(new_n605_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n604_), .A2(new_n572_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n255_), .A2(new_n248_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n702_), .A2(new_n248_), .B1(new_n707_), .B2(new_n708_), .ZN(G1332gat));
  OR3_X1    g508(.A1(new_n707_), .A2(G64gat), .A3(new_n602_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n700_), .A2(new_n701_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n427_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G64gat), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(KEYINPUT48), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(KEYINPUT48), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(G1333gat));
  OR3_X1    g515(.A1(new_n707_), .A2(G71gat), .A3(new_n634_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n701_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n388_), .A3(new_n699_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G71gat), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT114), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT114), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n722_), .A3(G71gat), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n721_), .A2(KEYINPUT49), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT49), .B1(new_n721_), .B2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n717_), .B1(new_n724_), .B2(new_n725_), .ZN(G1334gat));
  OR3_X1    g525(.A1(new_n707_), .A2(G78gat), .A3(new_n638_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n711_), .A2(new_n639_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G78gat), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT50), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT50), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1335gat));
  AND2_X1   g531(.A1(new_n543_), .A2(new_n544_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n733_), .A2(new_n572_), .A3(new_n589_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n655_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n433_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n705_), .A2(new_n609_), .A3(new_n645_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n250_), .A3(new_n255_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n736_), .B2(new_n602_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n326_), .A3(new_n427_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  NAND2_X1  g542(.A1(new_n735_), .A2(new_n388_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n634_), .A2(new_n436_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n744_), .A2(G99gat), .B1(new_n738_), .B2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT115), .B1(new_n746_), .B2(KEYINPUT116), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT51), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n746_), .B2(KEYINPUT115), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n747_), .B2(new_n750_), .ZN(G1338gat));
  INV_X1    g550(.A(new_n437_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n738_), .A2(new_n752_), .A3(new_n416_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n735_), .A2(new_n416_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G106gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n753_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  XOR2_X1   g561(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n763_));
  NAND2_X1  g562(.A1(new_n572_), .A2(new_n536_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n521_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n508_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n765_), .A2(KEYINPUT55), .B1(new_n766_), .B2(new_n511_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n522_), .A2(new_n768_), .A3(new_n527_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n534_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n534_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n764_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n556_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n555_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n568_), .C1(new_n776_), .C2(new_n562_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n571_), .A2(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n535_), .A2(KEYINPUT73), .A3(new_n536_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT73), .B1(new_n535_), .B2(new_n536_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT118), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n779_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n775_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n493_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n763_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n775_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n784_), .B1(new_n541_), .B2(new_n779_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n785_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n493_), .A2(KEYINPUT57), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT120), .B1(new_n786_), .B2(new_n794_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n773_), .A2(new_n774_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n779_), .A2(new_n536_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n798_), .A2(KEYINPUT58), .A3(new_n799_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n606_), .A3(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n788_), .A2(new_n796_), .A3(new_n797_), .A4(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n543_), .A2(new_n544_), .A3(new_n697_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT117), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n543_), .A2(new_n808_), .A3(new_n544_), .A4(new_n697_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n605_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT54), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n807_), .A2(new_n812_), .A3(new_n605_), .A4(new_n809_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n805_), .A2(new_n607_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n429_), .A2(new_n433_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n602_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT59), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n819_), .B2(new_n816_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n796_), .A2(new_n797_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n792_), .A2(new_n493_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n605_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n823_), .A2(new_n763_), .B1(new_n803_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n589_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n811_), .A2(new_n813_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n817_), .A2(new_n572_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G113gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n805_), .A2(new_n607_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n811_), .A2(new_n813_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n816_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OR3_X1    g634(.A1(new_n835_), .A2(G113gat), .A3(new_n610_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n830_), .A2(new_n836_), .ZN(G1340gat));
  NAND3_X1  g636(.A1(new_n817_), .A2(new_n609_), .A3(new_n828_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G120gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n733_), .A2(G120gat), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n840_), .B(G120gat), .S(KEYINPUT60), .Z(new_n841_));
  NAND3_X1  g640(.A1(new_n833_), .A2(new_n834_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n814_), .A2(new_n816_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(KEYINPUT122), .A3(new_n841_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n847_), .ZN(G1341gat));
  NAND3_X1  g647(.A1(new_n817_), .A2(new_n589_), .A3(new_n828_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G127gat), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n835_), .A2(G127gat), .A3(new_n607_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(new_n845_), .B2(new_n787_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n817_), .A2(new_n828_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT123), .B(G134gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n605_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n854_), .B2(new_n856_), .ZN(G1343gat));
  INV_X1    g656(.A(new_n431_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n602_), .A2(new_n255_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n833_), .A2(new_n572_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n833_), .A2(new_n609_), .A3(new_n860_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT124), .B(G148gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1345gat));
  NAND3_X1  g664(.A1(new_n833_), .A2(new_n589_), .A3(new_n860_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n833_), .A2(new_n869_), .A3(new_n787_), .A4(new_n860_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n814_), .A2(new_n605_), .A3(new_n859_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1347gat));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n602_), .A2(new_n255_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n388_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n639_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n814_), .A2(new_n610_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n878_), .B2(new_n266_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n833_), .A2(new_n876_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT62), .B(G169gat), .C1(new_n880_), .C2(new_n610_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n268_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  AOI21_X1  g682(.A(new_n877_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G176gat), .B1(new_n884_), .B2(new_n609_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n814_), .A2(new_n416_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n733_), .A2(new_n875_), .A3(new_n265_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  NOR3_X1   g687(.A1(new_n880_), .A2(new_n607_), .A3(new_n278_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n875_), .A2(new_n607_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G183gat), .B1(new_n886_), .B2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1350gat));
  NAND2_X1  g691(.A1(new_n787_), .A2(new_n279_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT126), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n884_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  INV_X1    g695(.A(G190gat), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n896_), .B(new_n897_), .C1(new_n884_), .C2(new_n606_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n606_), .B(new_n876_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT125), .B1(new_n899_), .B2(G190gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n895_), .B1(new_n898_), .B2(new_n900_), .ZN(G1351gat));
  NAND2_X1  g700(.A1(new_n874_), .A2(new_n858_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n833_), .A2(G197gat), .A3(new_n572_), .A4(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n814_), .A2(new_n902_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n907_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n572_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n833_), .A2(new_n572_), .A3(new_n903_), .ZN(new_n909_));
  INV_X1    g708(.A(G197gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n906_), .A2(new_n908_), .A3(new_n911_), .ZN(G1352gat));
  AND3_X1   g711(.A1(new_n907_), .A2(G204gat), .A3(new_n609_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G204gat), .B1(new_n907_), .B2(new_n609_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1353gat));
  OR2_X1    g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n907_), .B2(new_n589_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n907_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n607_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT63), .B(G211gat), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  OAI21_X1  g720(.A(G218gat), .B1(new_n918_), .B2(new_n605_), .ZN(new_n922_));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n907_), .A2(new_n923_), .A3(new_n787_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1355gat));
endmodule


