//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT101), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT89), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT2), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(KEYINPUT2), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n212_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n218_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .A4(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n208_), .B(new_n209_), .C1(new_n216_), .C2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n212_), .A2(new_n222_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT90), .ZN(new_n228_));
  AND3_X1   g027(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n208_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n227_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n226_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT93), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n226_), .B(KEYINPUT93), .C1(new_n233_), .C2(new_n232_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n207_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(KEYINPUT4), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n226_), .B(new_n207_), .C1(new_n233_), .C2(new_n232_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT4), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n204_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n238_), .A2(new_n203_), .A3(new_n241_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  INV_X1    g045(.A(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G57gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n207_), .B(KEYINPUT31), .Z(new_n255_));
  XNOR2_X1  g054(.A(G71gat), .B(G99gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G43gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT30), .B(G15gat), .Z(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT82), .B(G183gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT25), .ZN(new_n262_));
  OR2_X1    g061(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G190gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT83), .A3(KEYINPUT26), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(KEYINPUT26), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(KEYINPUT26), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT83), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .A4(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT84), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  INV_X1    g073(.A(G169gat), .ZN(new_n275_));
  INV_X1    g074(.A(G176gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(G169gat), .B2(G176gat), .ZN(new_n280_));
  INV_X1    g079(.A(G183gat), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n281_), .A2(new_n265_), .A3(KEYINPUT23), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT23), .B1(new_n281_), .B2(new_n265_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n280_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n273_), .A2(new_n274_), .A3(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n283_), .B(KEYINPUT85), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n282_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(G190gat), .B2(new_n261_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT22), .B(G169gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n277_), .B1(new_n291_), .B2(new_n276_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n287_), .A2(KEYINPUT86), .A3(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n260_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n287_), .A2(KEYINPUT86), .A3(new_n293_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT86), .B1(new_n287_), .B2(new_n293_), .ZN(new_n303_));
  OAI211_X1 g102(.A(G227gat), .B(G233gat), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n259_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(KEYINPUT87), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n255_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n301_), .A2(KEYINPUT88), .A3(new_n306_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(new_n312_), .B2(new_n255_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n236_), .A2(new_n314_), .A3(new_n237_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n236_), .A2(new_n314_), .A3(new_n237_), .A4(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G22gat), .B(G50gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(new_n321_), .A3(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n326_));
  AND2_X1   g125(.A1(new_n234_), .A2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G197gat), .B(G204gat), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT21), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n328_), .A2(KEYINPUT21), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n330_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(G228gat), .B(G233gat), .C1(new_n327_), .C2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G78gat), .B(G106gat), .Z(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT96), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n314_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n336_), .B(new_n339_), .C1(new_n340_), .C2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n336_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n337_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n325_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n338_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n343_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT97), .B1(new_n350_), .B2(new_n325_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n325_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT97), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n347_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n254_), .B1(new_n313_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT19), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT20), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n296_), .A2(new_n297_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(new_n334_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n267_), .A2(new_n268_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT25), .B(G183gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n289_), .A2(new_n280_), .A3(new_n285_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT98), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n292_), .B(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n284_), .B1(G183gat), .B2(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT102), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n334_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n372_), .B2(new_n371_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n359_), .B1(new_n362_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n360_), .B1(new_n371_), .B2(new_n334_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n361_), .B2(new_n334_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(new_n358_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380_));
  INV_X1    g179(.A(G92gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT18), .B(G64gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT103), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT103), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n387_), .B(new_n384_), .C1(new_n375_), .C2(new_n378_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n335_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT99), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n358_), .B1(new_n362_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n358_), .B(new_n376_), .C1(new_n361_), .C2(new_n334_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n388_), .A2(KEYINPUT27), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n302_), .A2(new_n303_), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT20), .B(new_n390_), .C1(new_n396_), .C2(new_n335_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n359_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n384_), .A3(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT100), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT100), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n398_), .A2(new_n401_), .A3(new_n384_), .A4(new_n392_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n402_), .A3(new_n394_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT27), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n386_), .A2(new_n395_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n354_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n353_), .B1(new_n352_), .B2(new_n349_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n255_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n410_));
  OAI22_X1  g209(.A1(new_n408_), .A2(new_n347_), .B1(new_n410_), .B2(new_n309_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n356_), .A2(new_n405_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n254_), .B(new_n414_), .C1(new_n379_), .C2(new_n413_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n252_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n245_), .A2(KEYINPUT33), .A3(new_n251_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n238_), .A2(new_n241_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n251_), .B1(new_n419_), .B2(new_n203_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n239_), .A2(new_n242_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n203_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n415_), .B1(new_n423_), .B2(new_n403_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n355_), .A3(new_n313_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n412_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT72), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT70), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n247_), .A2(new_n381_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G85gat), .A2(G92gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G99gat), .A2(G106gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n436_));
  NOR3_X1   g235(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT7), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n435_), .B(new_n436_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n437_), .A2(new_n438_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n432_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT64), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n429_), .A2(new_n444_), .A3(new_n430_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT9), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT9), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n429_), .A2(new_n444_), .A3(new_n447_), .A4(new_n430_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n429_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n435_), .A2(new_n436_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT10), .B(G99gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G106gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n450_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  OAI221_X1 g254(.A(new_n432_), .B1(KEYINPUT66), .B2(KEYINPUT8), .C1(new_n439_), .C2(new_n440_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n443_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT67), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT67), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n443_), .A2(new_n455_), .A3(new_n456_), .A4(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G57gat), .ZN(new_n462_));
  INV_X1    g261(.A(G64gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G57gat), .A2(G64gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G71gat), .B(G78gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT11), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n464_), .A2(new_n470_), .A3(new_n465_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT11), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT68), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(KEYINPUT68), .A3(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT69), .B1(new_n461_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481_));
  AOI211_X1 g280(.A(new_n481_), .B(new_n478_), .C1(new_n458_), .C2(new_n460_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n428_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n442_), .A2(new_n441_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n459_), .B1(new_n484_), .B2(new_n456_), .ZN(new_n485_));
  AND4_X1   g284(.A1(new_n459_), .A2(new_n443_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n479_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n481_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n461_), .A2(KEYINPUT69), .A3(new_n479_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT70), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n458_), .A2(new_n460_), .A3(new_n478_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(G230gat), .A2(G233gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n474_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n457_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n493_), .B1(new_n461_), .B2(new_n479_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n491_), .A2(KEYINPUT71), .A3(new_n495_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT71), .B1(new_n491_), .B2(new_n495_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n497_), .B(new_n498_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G120gat), .B(G148gat), .ZN(new_n502_));
  INV_X1    g301(.A(G204gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT5), .B(G176gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  AND4_X1   g305(.A1(new_n427_), .A2(new_n494_), .A3(new_n501_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n491_), .A2(new_n495_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n491_), .A2(KEYINPUT71), .A3(new_n495_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n510_), .A2(new_n511_), .B1(new_n457_), .B2(new_n496_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n492_), .A2(new_n493_), .B1(new_n512_), .B2(new_n498_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n427_), .B1(new_n513_), .B2(new_n506_), .ZN(new_n514_));
  OAI22_X1  g313(.A1(new_n507_), .A2(new_n514_), .B1(new_n513_), .B2(new_n506_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n516_));
  OR2_X1    g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT81), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(KEYINPUT76), .A2(G15gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT76), .A2(G15gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G22gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT77), .B(G8gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT14), .ZN(new_n529_));
  INV_X1    g328(.A(G22gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n530_), .A3(new_n525_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(G1gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(KEYINPUT14), .A2(G1gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n527_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(G8gat), .ZN(new_n537_));
  INV_X1    g336(.A(G8gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n538_), .A3(new_n535_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G29gat), .B(G36gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G43gat), .B(G50gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n523_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n542_), .B(KEYINPUT15), .ZN(new_n547_));
  INV_X1    g346(.A(new_n539_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n538_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(new_n543_), .A3(new_n522_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n521_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n537_), .A2(new_n539_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n542_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n522_), .B1(new_n555_), .B2(new_n543_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT80), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G169gat), .B(G197gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n552_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n551_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT80), .B1(new_n563_), .B2(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n546_), .A2(new_n521_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n520_), .B1(new_n561_), .B2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n560_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(new_n565_), .A3(new_n562_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(KEYINPUT81), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(G211gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT79), .B(G183gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n475_), .B1(new_n577_), .B2(KEYINPUT17), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(new_n553_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n553_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n474_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n581_), .A2(new_n473_), .A3(new_n472_), .A4(new_n582_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n461_), .A2(new_n542_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT35), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n547_), .A2(new_n457_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n594_), .A2(new_n590_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT36), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT75), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n598_), .A2(new_n607_), .A3(new_n599_), .A4(new_n603_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n605_), .A2(KEYINPUT75), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n588_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n605_), .A2(KEYINPUT37), .A3(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n587_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n426_), .A2(new_n519_), .A3(new_n571_), .A4(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT104), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT104), .ZN(new_n617_));
  INV_X1    g416(.A(new_n254_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(G1gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT105), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT105), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n519_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n571_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n609_), .A2(new_n610_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n587_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n426_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n618_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n621_), .A2(KEYINPUT38), .A3(new_n622_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n625_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n405_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(new_n528_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n616_), .A2(new_n617_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n616_), .A2(KEYINPUT106), .A3(new_n617_), .A4(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G8gat), .B1(new_n631_), .B2(new_n405_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT39), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n641_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1325gat));
  AND2_X1   g446(.A1(new_n616_), .A2(new_n617_), .ZN(new_n648_));
  INV_X1    g447(.A(G15gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n313_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n631_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n649_), .B1(new_n655_), .B2(new_n650_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n653_), .A2(new_n654_), .A3(new_n658_), .A4(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(new_n355_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n648_), .A2(new_n530_), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G22gat), .B1(new_n631_), .B2(new_n355_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(KEYINPUT42), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT42), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n426_), .A2(new_n613_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n426_), .A2(KEYINPUT43), .A3(new_n613_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(new_n628_), .A3(new_n587_), .A4(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n587_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n628_), .A4(new_n670_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n254_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G29gat), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n628_), .A2(new_n426_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n629_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n674_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n618_), .A2(G29gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  NAND3_X1  g483(.A1(new_n673_), .A2(new_n635_), .A3(new_n676_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n405_), .A2(G36gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n682_), .A2(KEYINPUT45), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT45), .B1(new_n682_), .B2(new_n688_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n686_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n686_), .A2(new_n691_), .A3(KEYINPUT46), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1329gat));
  NOR3_X1   g495(.A1(new_n682_), .A2(G43gat), .A3(new_n313_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n673_), .A2(new_n650_), .A3(new_n676_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(G43gat), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT47), .B(new_n697_), .C1(new_n698_), .C2(G43gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1330gat));
  NAND3_X1  g502(.A1(new_n673_), .A2(new_n661_), .A3(new_n676_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G50gat), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n355_), .A2(G50gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n682_), .B2(new_n706_), .ZN(G1331gat));
  AOI21_X1  g506(.A(new_n571_), .B1(new_n412_), .B2(new_n425_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT109), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n626_), .A3(new_n614_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n462_), .B1(new_n710_), .B2(new_n618_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n708_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(G57gat), .A3(new_n254_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n713_), .A2(new_n714_), .A3(new_n716_), .ZN(G1332gat));
  AOI21_X1  g516(.A(new_n463_), .B1(new_n715_), .B2(new_n635_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT48), .Z(new_n719_));
  NAND2_X1  g518(.A1(new_n635_), .A2(new_n463_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n710_), .B2(new_n720_), .ZN(G1333gat));
  INV_X1    g520(.A(G71gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n715_), .B2(new_n650_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT49), .Z(new_n724_));
  NAND2_X1  g523(.A1(new_n650_), .A2(new_n722_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n710_), .B2(new_n725_), .ZN(G1334gat));
  INV_X1    g525(.A(G78gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n715_), .B2(new_n661_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n661_), .A2(new_n727_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n710_), .B2(new_n731_), .ZN(G1335gat));
  NAND3_X1  g531(.A1(new_n709_), .A2(new_n626_), .A3(new_n681_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n254_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n626_), .A2(new_n627_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n669_), .A2(new_n587_), .A3(new_n670_), .A4(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n675_), .A2(KEYINPUT112), .A3(new_n670_), .A4(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n618_), .A2(new_n247_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n735_), .B1(new_n744_), .B2(new_n745_), .ZN(G1336gat));
  AOI21_X1  g545(.A(G92gat), .B1(new_n734_), .B2(new_n635_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n405_), .A2(new_n381_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n744_), .B2(new_n748_), .ZN(G1337gat));
  NAND3_X1  g548(.A1(new_n740_), .A2(new_n650_), .A3(new_n741_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G99gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n734_), .A2(new_n452_), .A3(new_n650_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT51), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n755_), .A3(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1338gat));
  NAND4_X1  g556(.A1(new_n675_), .A2(new_n661_), .A3(new_n670_), .A4(new_n737_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G106gat), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n661_), .A2(new_n453_), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n760_), .A2(new_n761_), .B1(new_n733_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI221_X1 g564(.A(new_n765_), .B1(new_n733_), .B2(new_n762_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  OAI221_X1 g567(.A(new_n497_), .B1(new_n480_), .B2(new_n482_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n493_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n501_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n510_), .A2(new_n511_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n497_), .A4(new_n498_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n770_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n768_), .A3(new_n493_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n506_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n497_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n480_), .A2(new_n482_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n493_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT115), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(new_n777_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n506_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT56), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n522_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n550_), .A2(new_n523_), .A3(new_n543_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n560_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n569_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n494_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT72), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n513_), .A2(new_n427_), .A3(new_n506_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n780_), .A2(new_n788_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n780_), .A2(new_n788_), .A3(KEYINPUT58), .A4(new_n796_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n613_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n779_), .B1(new_n778_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n571_), .B1(new_n507_), .B2(new_n514_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT114), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n571_), .B(new_n806_), .C1(new_n507_), .C2(new_n514_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n787_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n803_), .A2(new_n805_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n515_), .A2(new_n569_), .A3(new_n791_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n629_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n801_), .B1(new_n811_), .B2(KEYINPUT57), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n813_), .B(new_n629_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n587_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n614_), .A2(new_n627_), .A3(new_n519_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n614_), .A2(new_n818_), .A3(new_n627_), .A4(new_n519_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n635_), .A2(new_n618_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n821_), .A2(new_n355_), .A3(new_n650_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n661_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(new_n650_), .A3(new_n822_), .A4(new_n825_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n627_), .A2(new_n832_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n823_), .A2(new_n627_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n831_), .A2(new_n833_), .B1(new_n834_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836_));
  AOI21_X1  g635(.A(G120gat), .B1(new_n626_), .B2(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n837_), .A2(KEYINPUT118), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT60), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n837_), .A2(KEYINPUT118), .ZN(new_n841_));
  OR4_X1    g640(.A1(new_n823_), .A2(new_n838_), .A3(new_n840_), .A4(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n519_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n839_), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n587_), .A2(new_n845_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n823_), .A2(new_n587_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n831_), .A2(new_n846_), .B1(new_n847_), .B2(new_n845_), .ZN(G1342gat));
  INV_X1    g647(.A(new_n613_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT119), .B(G134gat), .Z(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n823_), .A2(new_n680_), .ZN(new_n852_));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n831_), .A2(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1343gat));
  NOR2_X1   g653(.A1(new_n650_), .A2(new_n355_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(new_n822_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n571_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n626_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g661(.A1(new_n821_), .A2(new_n674_), .A3(new_n822_), .A4(new_n855_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n857_), .A2(new_n865_), .A3(new_n674_), .A4(new_n822_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n864_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1346gat));
  AOI21_X1  g669(.A(G162gat), .B1(new_n858_), .B2(new_n629_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n613_), .A2(G162gat), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n858_), .B2(new_n872_), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n405_), .A2(new_n254_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n571_), .A3(new_n650_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n829_), .A2(new_n291_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(KEYINPUT121), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n875_), .A2(KEYINPUT121), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n829_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n880_), .A2(new_n881_), .A3(G169gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(G169gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n877_), .B1(new_n882_), .B2(new_n883_), .ZN(G1348gat));
  NAND4_X1  g683(.A1(new_n829_), .A2(new_n626_), .A3(new_n650_), .A4(new_n874_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT122), .B(G176gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1349gat));
  NAND4_X1  g686(.A1(new_n829_), .A2(new_n650_), .A3(new_n674_), .A4(new_n874_), .ZN(new_n888_));
  MUX2_X1   g687(.A(new_n364_), .B(new_n261_), .S(new_n888_), .Z(G1350gat));
  AND2_X1   g688(.A1(new_n829_), .A2(new_n650_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n890_), .A2(new_n363_), .A3(new_n629_), .A4(new_n874_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n890_), .A2(new_n613_), .A3(new_n874_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n265_), .ZN(G1351gat));
  INV_X1    g692(.A(new_n874_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n856_), .B(new_n894_), .C1(new_n815_), .C2(new_n820_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n571_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  XOR2_X1   g696(.A(KEYINPUT123), .B(G204gat), .Z(new_n898_));
  NAND2_X1  g697(.A1(new_n503_), .A2(KEYINPUT123), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n626_), .ZN(new_n900_));
  MUX2_X1   g699(.A(new_n898_), .B(new_n899_), .S(new_n900_), .Z(G1353gat));
  XOR2_X1   g700(.A(KEYINPUT63), .B(G211gat), .Z(new_n902_));
  NAND4_X1  g701(.A1(new_n857_), .A2(new_n674_), .A3(new_n874_), .A4(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT124), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n895_), .A2(new_n905_), .A3(new_n674_), .A4(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n821_), .A2(new_n674_), .A3(new_n855_), .A4(new_n874_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT125), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n908_), .A2(KEYINPUT125), .A3(new_n909_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n907_), .A2(new_n910_), .A3(new_n911_), .ZN(G1354gat));
  XOR2_X1   g711(.A(KEYINPUT127), .B(G218gat), .Z(new_n913_));
  AND3_X1   g712(.A1(new_n895_), .A2(new_n613_), .A3(new_n913_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n857_), .A2(new_n629_), .A3(new_n874_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n913_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n895_), .A2(new_n629_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n914_), .B1(new_n917_), .B2(new_n919_), .ZN(G1355gat));
endmodule


