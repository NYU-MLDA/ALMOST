//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_;
  AND3_X1   g000(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT82), .B1(G183gat), .B2(G190gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT83), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(new_n212_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n213_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  INV_X1    g026(.A(G176gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n215_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(KEYINPUT24), .A3(new_n220_), .A4(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n223_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n206_), .B1(new_n202_), .B2(new_n203_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n218_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  INV_X1    g037(.A(G43gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G127gat), .B(G134gat), .Z(new_n244_));
  XOR2_X1   g043(.A(G113gat), .B(G120gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(G15gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT30), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n247_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n243_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G22gat), .B(G50gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G228gat), .A2(G233gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G218gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G211gat), .ZN(new_n263_));
  INV_X1    g062(.A(G211gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G218gat), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268_));
  NOR4_X1   g067(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n270_));
  AND2_X1   g069(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n271_), .A2(new_n272_), .A3(G197gat), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT21), .B1(new_n258_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n266_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(G197gat), .B1(new_n271_), .B2(new_n272_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n268_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT21), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n270_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n267_), .B1(new_n261_), .B2(new_n268_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n263_), .A2(new_n265_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n259_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n267_), .B1(G197gat), .B2(G204gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(KEYINPUT90), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n269_), .B1(new_n280_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT86), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n289_), .A2(G155gat), .A3(G162gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(G155gat), .B2(G162gat), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n290_), .A2(new_n291_), .B1(G155gat), .B2(G162gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT3), .ZN(new_n293_));
  INV_X1    g092(.A(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G148gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT87), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n293_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT88), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n292_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n298_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n308_), .A2(new_n309_), .B1(G141gat), .B2(G148gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n290_), .A2(new_n291_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT1), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n288_), .B1(new_n306_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n257_), .B1(new_n287_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G78gat), .ZN(new_n317_));
  INV_X1    g116(.A(G78gat), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(new_n257_), .C1(new_n287_), .C2(new_n315_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n317_), .A2(G106gat), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(G106gat), .B1(new_n317_), .B2(new_n319_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n254_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n306_), .A2(new_n314_), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n323_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT28), .B1(new_n323_), .B2(KEYINPUT29), .ZN(new_n325_));
  NAND3_X1  g124(.A1(KEYINPUT91), .A2(G228gat), .A3(G233gat), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G106gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n323_), .A2(KEYINPUT29), .ZN(new_n331_));
  INV_X1    g130(.A(new_n269_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n276_), .A2(new_n279_), .A3(new_n270_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT90), .B1(new_n281_), .B2(new_n285_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n318_), .B1(new_n336_), .B2(new_n257_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n319_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n330_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n317_), .A2(G106gat), .A3(new_n319_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n254_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n322_), .A2(new_n329_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n329_), .B1(new_n322_), .B2(new_n342_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n323_), .A2(new_n247_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n306_), .A2(new_n246_), .A3(new_n314_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT4), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n323_), .A2(new_n348_), .A3(new_n247_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT95), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT96), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n345_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n343_), .A2(new_n344_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT20), .B1(new_n335_), .B2(new_n237_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n228_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n230_), .B(KEYINPUT93), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n205_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT23), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n234_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n209_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n371_), .B1(new_n377_), .B2(KEYINPUT94), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n208_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n382_));
  INV_X1    g181(.A(G183gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(KEYINPUT25), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(KEYINPUT25), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n225_), .A2(KEYINPUT92), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n224_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n219_), .A2(new_n215_), .A3(new_n228_), .ZN(new_n389_));
  AND4_X1   g188(.A1(new_n207_), .A2(new_n231_), .A3(new_n204_), .A4(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n378_), .A2(new_n381_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(new_n287_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n366_), .B1(new_n367_), .B2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G8gat), .B(G36gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT18), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n366_), .B1(new_n391_), .B2(new_n287_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n335_), .B2(new_n237_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(new_n397_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT27), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT98), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n287_), .B1(new_n391_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n390_), .A2(new_n388_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n369_), .B(new_n370_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n377_), .A2(KEYINPUT94), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n406_), .B(new_n404_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n400_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n216_), .B1(new_n210_), .B2(KEYINPUT83), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n412_), .A2(new_n213_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n399_), .B1(new_n287_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n366_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n335_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n411_), .A2(new_n366_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n414_), .A2(new_n417_), .A3(KEYINPUT99), .A4(new_n415_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n397_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n403_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT27), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n398_), .A2(new_n400_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n415_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n423_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n397_), .B1(new_n393_), .B2(new_n401_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n425_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT100), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n423_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n402_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT100), .A3(new_n425_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n424_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n364_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n397_), .A2(KEYINPUT32), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n393_), .A2(new_n438_), .A3(new_n401_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n359_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n345_), .A2(new_n346_), .A3(new_n352_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n358_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT97), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n347_), .A2(new_n351_), .A3(new_n349_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT97), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n353_), .A2(KEYINPUT33), .A3(new_n354_), .A4(new_n358_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n443_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  OAI22_X1  g252(.A1(new_n439_), .A2(new_n441_), .B1(new_n453_), .B2(new_n434_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n253_), .B1(new_n437_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT100), .B1(new_n434_), .B2(new_n425_), .ZN(new_n457_));
  AOI211_X1 g256(.A(new_n431_), .B(KEYINPUT27), .C1(new_n433_), .C2(new_n402_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n397_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n459_));
  OAI22_X1  g258(.A1(new_n457_), .A2(new_n458_), .B1(new_n459_), .B2(new_n403_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n343_), .A2(new_n344_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n253_), .A2(new_n362_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n456_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G15gat), .B(G22gat), .ZN(new_n471_));
  INV_X1    g270(.A(G1gat), .ZN(new_n472_));
  INV_X1    g271(.A(G8gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G8gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n470_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(new_n477_), .B2(new_n467_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n467_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n477_), .A2(new_n467_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n479_), .A2(new_n482_), .B1(new_n486_), .B2(new_n481_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G113gat), .B(G141gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(G169gat), .B(G197gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n487_), .B(new_n490_), .Z(new_n491_));
  NOR2_X1   g290(.A1(new_n464_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n494_));
  XOR2_X1   g293(.A(G71gat), .B(G78gat), .Z(new_n495_));
  OR2_X1    g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n495_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT78), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(new_n478_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G127gat), .B(G155gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT16), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G183gat), .B(G211gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT17), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT79), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n503_), .A2(KEYINPUT80), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512_));
  OR3_X1    g311(.A1(new_n503_), .A2(new_n512_), .A3(new_n507_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT80), .B1(new_n503_), .B2(new_n509_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n511_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G190gat), .B(G218gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G134gat), .B(G162gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT75), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT10), .B(G99gat), .Z(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT64), .B(G106gat), .Z(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(G99gat), .A3(G106gat), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n526_), .A2(new_n527_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533_));
  INV_X1    g332(.A(G85gat), .ZN(new_n534_));
  INV_X1    g333(.A(G92gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n536_), .B2(KEYINPUT9), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(KEYINPUT66), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G92gat), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n534_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n532_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n532_), .B2(new_n543_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G99gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n330_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT67), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n548_), .A2(new_n330_), .A3(KEYINPUT67), .A4(KEYINPUT7), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n529_), .A2(new_n531_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT8), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G85gat), .B(G92gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n555_), .A2(new_n554_), .B1(new_n557_), .B2(KEYINPUT68), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n529_), .A2(new_n531_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n560_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n562_), .B1(new_n566_), .B2(new_n559_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n547_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n470_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT74), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n525_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n469_), .B1(new_n547_), .B2(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n532_), .A2(new_n543_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n557_), .A2(KEYINPUT68), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n556_), .A2(new_n574_), .A3(new_n565_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n559_), .B1(new_n575_), .B2(new_n561_), .ZN(new_n576_));
  AOI211_X1 g375(.A(KEYINPUT8), .B(new_n560_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n573_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT69), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT69), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n573_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n572_), .B1(new_n582_), .B2(new_n467_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n571_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n483_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n587_));
  NOR4_X1   g386(.A1(new_n587_), .A2(new_n570_), .A3(new_n572_), .A4(new_n525_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n521_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n580_), .B1(new_n567_), .B2(new_n573_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n581_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n467_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n569_), .A3(new_n585_), .ZN(new_n594_));
  OAI211_X1 g393(.A(KEYINPUT35), .B(new_n524_), .C1(new_n572_), .C2(KEYINPUT74), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n583_), .A2(new_n571_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n518_), .B(KEYINPUT36), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n589_), .A2(new_n590_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n598_), .B(KEYINPUT76), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n596_), .A2(new_n597_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n590_), .B1(new_n589_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT77), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n596_), .A2(new_n597_), .A3(new_n601_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n521_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT37), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n589_), .A2(new_n590_), .A3(new_n599_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n515_), .B1(new_n604_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n499_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT12), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n582_), .A2(new_n499_), .B1(new_n568_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n582_), .B2(new_n499_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT71), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n582_), .A2(new_n499_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n614_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n624_));
  OAI211_X1 g423(.A(G230gat), .B(G233gat), .C1(new_n623_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT71), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n617_), .A2(new_n619_), .A3(new_n626_), .A4(new_n620_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT5), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n630_), .B(new_n631_), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n622_), .A2(new_n625_), .A3(new_n627_), .A4(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT13), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n613_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n492_), .A2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(G1gat), .A3(new_n362_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT38), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT38), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n636_), .B(KEYINPUT13), .ZN(new_n644_));
  INV_X1    g443(.A(new_n491_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n515_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n589_), .A2(new_n599_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT101), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n464_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n362_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n642_), .A2(new_n643_), .A3(new_n653_), .ZN(G1324gat));
  INV_X1    g453(.A(new_n640_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n473_), .A3(new_n460_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n460_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G8gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT39), .B(new_n473_), .C1(new_n651_), .C2(new_n460_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g461(.A(new_n253_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G15gat), .B1(new_n652_), .B2(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT102), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT102), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(KEYINPUT41), .A3(new_n666_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n655_), .A2(new_n249_), .A3(new_n253_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n461_), .B(KEYINPUT103), .Z(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n651_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT42), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n655_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n513_), .A2(new_n514_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n510_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n646_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  INV_X1    g482(.A(new_n344_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n322_), .A2(new_n342_), .A3(new_n329_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n362_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n455_), .B1(new_n686_), .B2(new_n460_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n663_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n463_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n600_), .A2(new_n603_), .A3(KEYINPUT77), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n609_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n604_), .A2(KEYINPUT105), .A3(new_n611_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n690_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n688_), .A2(new_n689_), .A3(KEYINPUT104), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n683_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n604_), .A2(new_n611_), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT43), .B(new_n700_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT44), .B(new_n682_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n604_), .A2(KEYINPUT105), .A3(new_n611_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT105), .B1(new_n604_), .B2(new_n611_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n456_), .B2(new_n463_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n708_), .A3(new_n698_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n701_), .B1(new_n709_), .B2(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(new_n682_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n703_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n702_), .A2(new_n712_), .A3(G29gat), .A4(new_n363_), .ZN(new_n713_));
  INV_X1    g512(.A(G29gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n648_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n515_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n638_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n492_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n718_), .B2(new_n362_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n713_), .A2(new_n719_), .ZN(G1328gat));
  NAND3_X1  g519(.A1(new_n702_), .A2(new_n712_), .A3(new_n460_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G36gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n436_), .A2(G36gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n492_), .A2(new_n717_), .A3(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT45), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(KEYINPUT106), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(KEYINPUT106), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT107), .Z(new_n731_));
  NAND3_X1  g530(.A1(new_n726_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n731_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n725_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n721_), .B2(G36gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n735_), .B2(new_n728_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n736_), .ZN(G1329gat));
  NAND4_X1  g536(.A1(new_n702_), .A2(new_n712_), .A3(G43gat), .A4(new_n253_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n239_), .B1(new_n718_), .B2(new_n663_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1330gat));
  NAND4_X1  g541(.A1(new_n702_), .A2(new_n712_), .A3(G50gat), .A4(new_n461_), .ZN(new_n743_));
  INV_X1    g542(.A(G50gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n718_), .B2(new_n674_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1331gat));
  NOR4_X1   g545(.A1(new_n464_), .A2(new_n613_), .A3(new_n644_), .A4(new_n645_), .ZN(new_n747_));
  INV_X1    g546(.A(G57gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n363_), .ZN(new_n749_));
  AND4_X1   g548(.A1(new_n491_), .A2(new_n650_), .A3(new_n638_), .A4(new_n681_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n363_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n751_), .B2(new_n748_), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n750_), .B2(new_n460_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n747_), .A2(new_n753_), .A3(new_n460_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n750_), .B2(new_n253_), .ZN(new_n760_));
  XOR2_X1   g559(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n747_), .A2(new_n759_), .A3(new_n253_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1334gat));
  AOI21_X1  g563(.A(new_n318_), .B1(new_n750_), .B2(new_n675_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT50), .Z(new_n766_));
  NAND2_X1  g565(.A1(new_n675_), .A2(new_n318_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT111), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n747_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n644_), .A2(new_n716_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n688_), .A2(new_n689_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n491_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G85gat), .B1(new_n777_), .B2(new_n363_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n681_), .A2(new_n645_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n638_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n710_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n362_), .A2(new_n534_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT114), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n778_), .B1(new_n783_), .B2(new_n785_), .ZN(G1336gat));
  AOI21_X1  g585(.A(G92gat), .B1(new_n777_), .B2(new_n460_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n436_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n783_), .B2(new_n788_), .ZN(G1337gat));
  AND2_X1   g588(.A1(new_n253_), .A2(new_n526_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n777_), .A2(new_n790_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n710_), .A2(new_n782_), .A3(new_n663_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n548_), .ZN(new_n793_));
  OR2_X1    g592(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1338gat));
  NAND2_X1  g594(.A1(new_n461_), .A2(new_n527_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n461_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n710_), .A2(new_n782_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n799_), .B2(new_n330_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n780_), .B(KEYINPUT113), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n461_), .B(new_n801_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(G106gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n797_), .B1(new_n800_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n806_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n797_), .B(new_n808_), .C1(new_n800_), .C2(new_n804_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1339gat));
  NAND3_X1  g609(.A1(new_n644_), .A2(new_n612_), .A3(new_n491_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT118), .B1(new_n811_), .B2(KEYINPUT54), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n644_), .A2(new_n612_), .A3(new_n816_), .A4(new_n491_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n818_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n621_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n620_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n622_), .A2(new_n822_), .A3(new_n627_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n632_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n635_), .A2(KEYINPUT119), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n634_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT119), .A3(new_n829_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n645_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n490_), .B1(new_n486_), .B2(new_n480_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n479_), .A2(new_n485_), .A3(new_n481_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n487_), .A2(new_n490_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n636_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n715_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT57), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n491_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n842_), .A2(new_n833_), .B1(new_n636_), .B2(new_n837_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n715_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n832_), .A2(new_n829_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n635_), .A2(new_n837_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n832_), .B2(new_n829_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n700_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT58), .A3(new_n846_), .A4(new_n848_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n840_), .A2(new_n844_), .A3(new_n854_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n815_), .A2(new_n821_), .B1(new_n515_), .B2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n798_), .A2(new_n363_), .A3(new_n436_), .A4(new_n253_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(KEYINPUT59), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n843_), .A2(new_n841_), .A3(new_n715_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n854_), .B1(new_n839_), .B2(KEYINPUT57), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(KEYINPUT120), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n844_), .A2(new_n863_), .A3(new_n854_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n681_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n817_), .A2(new_n818_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n817_), .A2(new_n818_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n811_), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n868_), .B2(new_n812_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n859_), .B1(new_n865_), .B2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n858_), .A2(new_n871_), .A3(new_n645_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G113gat), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n856_), .A2(new_n857_), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n645_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(G1340gat));
  NAND3_X1  g676(.A1(new_n858_), .A2(new_n871_), .A3(new_n638_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G120gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n880_), .B2(G120gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(G120gat), .B1(new_n638_), .B2(new_n880_), .ZN(new_n882_));
  MUX2_X1   g681(.A(new_n881_), .B(KEYINPUT121), .S(new_n882_), .Z(new_n883_));
  NAND2_X1  g682(.A1(new_n874_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n884_), .ZN(G1341gat));
  NAND3_X1  g684(.A1(new_n858_), .A2(new_n871_), .A3(new_n681_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G127gat), .ZN(new_n887_));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n874_), .A2(new_n888_), .A3(new_n681_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n874_), .B2(new_n649_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n858_), .A2(new_n871_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT122), .B(G134gat), .Z(new_n893_));
  NOR2_X1   g692(.A1(new_n700_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n892_), .B2(new_n894_), .ZN(G1343gat));
  NOR4_X1   g694(.A1(new_n798_), .A2(new_n460_), .A3(new_n362_), .A4(new_n253_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT123), .Z(new_n897_));
  NAND2_X1  g696(.A1(new_n855_), .A2(new_n515_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n869_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n645_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT124), .B(G141gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n638_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n899_), .B2(new_n681_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n899_), .A2(new_n905_), .A3(new_n681_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n909_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n856_), .A2(KEYINPUT125), .A3(new_n515_), .A4(new_n897_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n906_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(G1346gat));
  AOI21_X1  g713(.A(G162gat), .B1(new_n899_), .B2(new_n649_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n706_), .A2(G162gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n899_), .B2(new_n916_), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n436_), .A2(new_n462_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n674_), .A2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n645_), .B(new_n919_), .C1(new_n865_), .C2(new_n870_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G169gat), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n865_), .A2(new_n870_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n924_), .A2(new_n368_), .A3(new_n645_), .A4(new_n919_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n920_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n923_), .A2(new_n925_), .A3(new_n926_), .ZN(G1348gat));
  NAND2_X1  g726(.A1(new_n869_), .A2(new_n898_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n928_), .A2(new_n798_), .A3(new_n918_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n929_), .A2(new_n228_), .A3(new_n644_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n924_), .A2(new_n638_), .A3(new_n919_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n228_), .B2(new_n931_), .ZN(G1349gat));
  AND2_X1   g731(.A1(new_n924_), .A2(new_n919_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n515_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n928_), .A2(new_n798_), .A3(new_n681_), .A4(new_n918_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n934_), .B1(new_n383_), .B2(new_n935_), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n924_), .A2(new_n851_), .A3(new_n919_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G190gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n649_), .A2(new_n224_), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(KEYINPUT126), .Z(new_n940_));
  NAND3_X1  g739(.A1(new_n924_), .A2(new_n919_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n686_), .A2(new_n436_), .A3(new_n253_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n869_), .B2(new_n898_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n645_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n638_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n949_), .B1(new_n274_), .B2(new_n948_), .ZN(G1353gat));
  NAND2_X1  g749(.A1(new_n945_), .A2(new_n681_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AND2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  AND2_X1   g754(.A1(new_n649_), .A2(new_n262_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n945_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n262_), .B1(new_n945_), .B2(new_n851_), .ZN(new_n959_));
  OAI21_X1  g758(.A(KEYINPUT127), .B1(new_n958_), .B2(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n856_), .A2(new_n700_), .A3(new_n944_), .ZN(new_n962_));
  OAI211_X1 g761(.A(new_n961_), .B(new_n957_), .C1(new_n962_), .C2(new_n262_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n960_), .A2(new_n963_), .ZN(G1355gat));
endmodule


