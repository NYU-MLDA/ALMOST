//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_;
  NOR2_X1   g000(.A1(G197gat), .A2(G204gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT88), .B(G204gat), .Z(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  NOR3_X1   g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(G169gat), .B2(G176gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G169gat), .B2(G176gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n211_), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT23), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n213_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(G183gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n223_), .B(new_n226_), .C1(new_n227_), .C2(new_n224_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(KEYINPUT80), .A3(new_n220_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n230_), .B(KEYINPUT23), .C1(new_n216_), .C2(new_n217_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n229_), .B(new_n231_), .C1(G183gat), .C2(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n239_));
  INV_X1    g038(.A(G169gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT22), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n234_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n222_), .A2(new_n228_), .B1(new_n232_), .B2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT89), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n205_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n205_), .A2(G204gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(G197gat), .B1(new_n244_), .B2(new_n245_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n247_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT21), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n208_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT90), .B1(new_n206_), .B2(new_n207_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n202_), .B1(new_n246_), .B2(G197gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT21), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n210_), .B(new_n243_), .C1(new_n254_), .C2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT20), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT94), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT93), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n208_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT89), .B1(new_n204_), .B2(G197gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n271_), .B2(KEYINPUT21), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n206_), .A2(KEYINPUT90), .A3(new_n207_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n257_), .B1(new_n256_), .B2(KEYINPUT21), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n209_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n229_), .A2(new_n231_), .A3(new_n215_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT96), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n229_), .A2(KEYINPUT96), .A3(new_n231_), .A4(new_n215_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n212_), .A2(KEYINPUT95), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(new_n214_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n212_), .A2(KEYINPUT95), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n283_), .A2(new_n284_), .B1(new_n227_), .B2(new_n223_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT22), .B(G169gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n234_), .B1(new_n287_), .B2(new_n237_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n281_), .A2(new_n285_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n276_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n260_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n263_), .A2(new_n268_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT20), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n276_), .B2(new_n289_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n210_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n243_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n267_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT18), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n291_), .A2(new_n292_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n294_), .B1(new_n276_), .B2(new_n243_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT94), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n267_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n305_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n295_), .A2(new_n268_), .A3(new_n298_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(KEYINPUT27), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT97), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n312_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n263_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(new_n267_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(KEYINPUT97), .A3(new_n311_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n290_), .B1(new_n308_), .B2(KEYINPUT94), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n268_), .B1(new_n322_), .B2(new_n263_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n305_), .B1(new_n323_), .B2(new_n318_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT27), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n315_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT84), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331_));
  INV_X1    g130(.A(G141gat), .ZN(new_n332_));
  INV_X1    g131(.A(G148gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(KEYINPUT83), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(KEYINPUT83), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n333_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n337_), .A2(KEYINPUT3), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n330_), .A2(new_n335_), .A3(new_n336_), .A4(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(G155gat), .B2(G162gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT1), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n339_), .B(new_n337_), .C1(new_n345_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT85), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT87), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n352_), .A2(KEYINPUT29), .A3(new_n354_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n363_), .B2(new_n296_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT91), .ZN(new_n366_));
  INV_X1    g165(.A(new_n351_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n296_), .B(new_n362_), .C1(new_n356_), .C2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT91), .B1(new_n370_), .B2(new_n364_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n359_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G22gat), .B(G50gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND3_X1  g175(.A1(new_n369_), .A2(new_n359_), .A3(new_n371_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n372_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G127gat), .B(G134gat), .Z(new_n383_));
  XOR2_X1   g182(.A(G113gat), .B(G120gat), .Z(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  NAND3_X1  g184(.A1(new_n352_), .A2(new_n354_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n367_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n352_), .A2(new_n392_), .A3(new_n354_), .A4(new_n385_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n386_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n394_), .A2(new_n395_), .A3(new_n400_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT100), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT100), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n406_), .A3(new_n403_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n385_), .B(KEYINPUT31), .Z(new_n409_));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410_));
  INV_X1    g209(.A(G43gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n243_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(G15gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n417_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n409_), .B1(new_n420_), .B2(KEYINPUT81), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(KEYINPUT81), .B2(new_n420_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n418_), .A2(new_n423_), .A3(new_n419_), .A4(new_n409_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n327_), .A2(new_n382_), .A3(new_n408_), .A4(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n311_), .A2(KEYINPUT32), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n402_), .A2(new_n403_), .B1(new_n301_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n427_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT98), .B1(new_n320_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT98), .ZN(new_n431_));
  NOR4_X1   g230(.A1(new_n323_), .A2(new_n431_), .A3(new_n318_), .A4(new_n427_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT99), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n403_), .A2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n394_), .A2(KEYINPUT33), .A3(new_n395_), .A4(new_n400_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n386_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n401_), .A3(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n436_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n441_), .A2(new_n321_), .A3(new_n324_), .A4(new_n317_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT99), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n428_), .B(new_n443_), .C1(new_n430_), .C2(new_n432_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n434_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  AND4_X1   g244(.A1(new_n378_), .A2(new_n381_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n445_), .A2(new_n382_), .B1(new_n446_), .B2(new_n327_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n426_), .B1(new_n447_), .B2(new_n425_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G29gat), .B(G36gat), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT71), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(KEYINPUT71), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G43gat), .B(G50gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460_));
  INV_X1    g259(.A(G1gat), .ZN(new_n461_));
  INV_X1    g260(.A(G8gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(KEYINPUT76), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT76), .ZN(new_n468_));
  INV_X1    g267(.A(new_n466_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(new_n458_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n458_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n449_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n456_), .A2(KEYINPUT15), .A3(new_n457_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT15), .B1(new_n456_), .B2(new_n457_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT77), .B1(new_n477_), .B2(new_n469_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT77), .B(new_n469_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n473_), .B1(new_n481_), .B2(new_n449_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G113gat), .B(G141gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n482_), .B(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n448_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT5), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G176gat), .B(G204gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT64), .B(G92gat), .Z(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT9), .B1(new_n493_), .B2(G85gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT9), .ZN(new_n495_));
  INV_X1    g294(.A(G85gat), .ZN(new_n496_));
  INV_X1    g295(.A(G92gat), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT65), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n498_), .B1(KEYINPUT65), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT6), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT10), .B(G99gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(G106gat), .B2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G85gat), .B(G92gat), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(G106gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT67), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(KEYINPUT66), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT7), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n521_), .B2(KEYINPUT67), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n517_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  AOI211_X1 g322(.A(KEYINPUT8), .B(new_n512_), .C1(new_n507_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(KEYINPUT68), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n517_), .B(new_n528_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n507_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n512_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT69), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n525_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n506_), .B1(new_n523_), .B2(KEYINPUT68), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n512_), .B1(new_n535_), .B2(new_n529_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n536_), .A2(KEYINPUT69), .A3(new_n526_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n511_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n538_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n545_), .B(new_n511_), .C1(new_n534_), .C2(new_n537_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(KEYINPUT70), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n538_), .A2(new_n552_), .A3(new_n546_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n548_), .A2(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n532_), .A2(new_n533_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT69), .B1(new_n536_), .B2(new_n526_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n525_), .A3(new_n557_), .ZN(new_n558_));
  AOI211_X1 g357(.A(KEYINPUT12), .B(new_n545_), .C1(new_n558_), .C2(new_n511_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n538_), .B2(new_n546_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n492_), .B1(new_n554_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n554_), .A2(new_n562_), .A3(new_n492_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT13), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(KEYINPUT36), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n530_), .A2(new_n531_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT8), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n524_), .B1(new_n573_), .B2(KEYINPUT69), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n510_), .B1(new_n574_), .B2(new_n556_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n459_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT35), .Z(new_n579_));
  INV_X1    g378(.A(KEYINPUT72), .ZN(new_n580_));
  AOI211_X1 g379(.A(new_n580_), .B(new_n476_), .C1(new_n558_), .C2(new_n511_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT72), .B1(new_n538_), .B2(new_n477_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n576_), .B(new_n579_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n538_), .A2(new_n458_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n575_), .B2(new_n476_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n538_), .A2(KEYINPUT72), .A3(new_n477_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n578_), .A2(KEYINPUT35), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n571_), .B(new_n583_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT73), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n576_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(KEYINPUT35), .A3(new_n578_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT73), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n571_), .A4(new_n583_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n570_), .B(KEYINPUT36), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n592_), .B2(new_n583_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n466_), .B(new_n545_), .Z(new_n605_));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT17), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n607_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n612_), .B(KEYINPUT17), .Z(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n607_), .B2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n598_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n604_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n487_), .A2(new_n567_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n408_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n461_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n448_), .A2(new_n600_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n567_), .A2(new_n486_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n616_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n408_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n622_), .A2(new_n623_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n624_), .A2(new_n630_), .A3(new_n631_), .ZN(G1324gat));
  NAND2_X1  g431(.A1(new_n325_), .A2(new_n326_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n314_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n628_), .A2(new_n448_), .A3(new_n634_), .A4(new_n600_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT101), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G8gat), .B1(new_n635_), .B2(KEYINPUT101), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT39), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n635_), .A2(KEYINPUT101), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(G8gat), .A4(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n620_), .A2(new_n462_), .A3(new_n634_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(KEYINPUT40), .A3(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1325gat));
  INV_X1    g448(.A(new_n425_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G15gat), .B1(new_n629_), .B2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT41), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n620_), .A2(new_n415_), .A3(new_n425_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  OAI21_X1  g453(.A(G22gat), .B1(new_n629_), .B2(new_n382_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT42), .ZN(new_n656_));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n382_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n620_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(G1327gat));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n626_), .A2(new_n616_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n604_), .A2(new_n618_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n448_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n448_), .B2(new_n664_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n662_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n621_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G29gat), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT13), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n566_), .B(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n617_), .A2(new_n627_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n487_), .A2(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(G29gat), .A3(new_n408_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n661_), .B1(new_n672_), .B2(new_n679_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT102), .B(new_n678_), .C1(new_n671_), .C2(G29gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1328gat));
  XNOR2_X1  g481(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n669_), .A2(new_n634_), .A3(new_n670_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n327_), .A2(G36gat), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n448_), .A2(new_n676_), .A3(new_n486_), .A4(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT45), .Z(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n683_), .B1(new_n685_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n683_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n688_), .B(new_n691_), .C1(new_n684_), .C2(G36gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1329gat));
  NAND4_X1  g492(.A1(new_n669_), .A2(G43gat), .A3(new_n425_), .A4(new_n670_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n411_), .B1(new_n677_), .B2(new_n650_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g496(.A1(new_n677_), .A2(new_n382_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(G50gat), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n669_), .A2(new_n670_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n658_), .A2(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(G1331gat));
  NOR3_X1   g501(.A1(new_n567_), .A2(new_n486_), .A3(new_n627_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n625_), .A2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT106), .B(G57gat), .Z(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n408_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(G57gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n486_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n448_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT104), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n674_), .A3(new_n619_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n711_), .B2(new_n408_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT105), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n707_), .C1(new_n711_), .C2(new_n408_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n706_), .B1(new_n713_), .B2(new_n715_), .ZN(G1332gat));
  OAI21_X1  g515(.A(G64gat), .B1(new_n704_), .B2(new_n327_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT48), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n327_), .A2(G64gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n711_), .B2(new_n719_), .ZN(G1333gat));
  OR3_X1    g519(.A1(new_n711_), .A2(G71gat), .A3(new_n650_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n625_), .A2(new_n425_), .A3(new_n703_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G71gat), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n723_), .A2(KEYINPUT108), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(KEYINPUT108), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n721_), .B1(new_n727_), .B2(new_n728_), .ZN(G1334gat));
  NAND3_X1  g528(.A1(new_n625_), .A2(new_n658_), .A3(new_n703_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G78gat), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT109), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT109), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n711_), .A2(G78gat), .A3(new_n382_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(KEYINPUT50), .A3(new_n733_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(G1335gat));
  OR2_X1    g538(.A1(new_n665_), .A2(new_n666_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n674_), .A2(new_n708_), .A3(new_n627_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT110), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n408_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n567_), .A2(new_n675_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n710_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n621_), .A2(new_n496_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(G1336gat));
  INV_X1    g547(.A(new_n743_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n634_), .A2(new_n493_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT111), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n710_), .A2(new_n634_), .A3(new_n745_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n749_), .A2(new_n751_), .B1(new_n752_), .B2(new_n497_), .ZN(G1337gat));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(KEYINPUT112), .ZN(new_n755_));
  OAI21_X1  g554(.A(G99gat), .B1(new_n743_), .B2(new_n650_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n650_), .A2(new_n508_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n746_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n755_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n756_), .B(new_n762_), .C1(new_n746_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1338gat));
  NAND4_X1  g563(.A1(new_n710_), .A2(new_n514_), .A3(new_n658_), .A4(new_n745_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n742_), .B(new_n658_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n765_), .B(new_n772_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n617_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n565_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n708_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n548_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n551_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n562_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n555_), .B(KEYINPUT55), .C1(new_n559_), .C2(new_n561_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT114), .B1(new_n786_), .B2(KEYINPUT113), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n785_), .A2(new_n491_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(KEYINPUT113), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n785_), .B2(new_n491_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n491_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT114), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n779_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n481_), .A2(KEYINPUT115), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n795_), .A2(G229gat), .A3(G233gat), .A4(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n471_), .A2(new_n472_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n485_), .B1(new_n799_), .B2(new_n449_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n798_), .A2(new_n800_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n777_), .B2(new_n563_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT116), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n566_), .A2(new_n804_), .A3(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n776_), .B1(new_n794_), .B2(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n801_), .A2(new_n565_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n491_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n491_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT58), .B(new_n808_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n603_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n617_), .A2(new_n601_), .A3(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n617_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n813_), .B(new_n814_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n785_), .A2(new_n491_), .A3(new_n787_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n782_), .A2(new_n562_), .B1(new_n780_), .B2(new_n551_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n492_), .B1(new_n820_), .B2(new_n784_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(new_n789_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n821_), .B2(KEYINPUT56), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n778_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n806_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n617_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n807_), .B(new_n818_), .C1(new_n827_), .C2(KEYINPUT57), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n619_), .A2(new_n829_), .A3(new_n708_), .A4(new_n567_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n604_), .A2(new_n567_), .A3(new_n616_), .A4(new_n618_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT54), .B1(new_n831_), .B2(new_n486_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n828_), .A2(new_n627_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n621_), .A2(new_n327_), .A3(new_n382_), .A4(new_n425_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT117), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n486_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n785_), .A2(new_n491_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n786_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n792_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT58), .B1(new_n844_), .B2(new_n808_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n814_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n825_), .A2(new_n826_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n847_), .A2(new_n664_), .B1(new_n848_), .B2(new_n776_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n794_), .A2(new_n806_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n775_), .B1(new_n850_), .B2(new_n617_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n616_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n830_), .A2(new_n832_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT59), .B(new_n835_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n708_), .B1(new_n841_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n839_), .B1(new_n855_), .B2(new_n838_), .ZN(G1340gat));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n567_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n837_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n857_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n567_), .B1(new_n841_), .B2(new_n854_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n837_), .A2(new_n862_), .A3(new_n616_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n627_), .B1(new_n841_), .B2(new_n854_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1342gat));
  NAND2_X1  g664(.A1(new_n664_), .A2(G134gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT118), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n807_), .A2(new_n818_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n848_), .B2(new_n600_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n627_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n830_), .A2(new_n832_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT59), .B1(new_n872_), .B2(new_n835_), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n840_), .B(new_n836_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n867_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876_));
  INV_X1    g675(.A(G134gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n835_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n600_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n876_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n867_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n841_), .B2(new_n854_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G134gat), .B1(new_n837_), .B2(new_n617_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT119), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n880_), .A2(new_n884_), .ZN(G1343gat));
  NOR4_X1   g684(.A1(new_n634_), .A2(new_n382_), .A3(new_n408_), .A4(new_n425_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT120), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n833_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n486_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n674_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT121), .B(G148gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n888_), .A2(new_n616_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(new_n887_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n872_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n664_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G162gat), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(G162gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n617_), .A2(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n900_), .B(KEYINPUT122), .C1(new_n898_), .C2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n888_), .B2(new_n664_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n898_), .A2(new_n902_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(G1347gat));
  XOR2_X1   g707(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n909_));
  NOR3_X1   g708(.A1(new_n327_), .A2(new_n621_), .A3(new_n650_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n382_), .B1(new_n910_), .B2(KEYINPUT123), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(KEYINPUT123), .B2(new_n910_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n872_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n708_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n909_), .B1(new_n914_), .B2(new_n240_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n287_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n909_), .ZN(new_n917_));
  OAI211_X1 g716(.A(G169gat), .B(new_n917_), .C1(new_n913_), .C2(new_n708_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n915_), .A2(new_n916_), .A3(new_n918_), .ZN(G1348gat));
  NOR2_X1   g718(.A1(new_n913_), .A2(new_n567_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n237_), .ZN(G1349gat));
  NOR3_X1   g720(.A1(new_n913_), .A2(new_n227_), .A3(new_n627_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n913_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n616_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n216_), .B2(new_n924_), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n223_), .A3(new_n617_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n872_), .A2(new_n664_), .A3(new_n912_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n927_), .A2(new_n928_), .A3(G190gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(G190gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n926_), .B1(new_n929_), .B2(new_n930_), .ZN(G1351gat));
  NAND3_X1  g730(.A1(new_n446_), .A2(new_n634_), .A3(new_n650_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n872_), .A2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n205_), .B1(new_n934_), .B2(new_n708_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n833_), .A2(new_n932_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n936_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n486_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(G197gat), .A3(new_n486_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(G1352gat));
  AND4_X1   g740(.A1(KEYINPUT127), .A2(new_n936_), .A3(new_n204_), .A4(new_n674_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n934_), .A2(new_n567_), .ZN(new_n943_));
  AOI21_X1  g742(.A(KEYINPUT127), .B1(new_n943_), .B2(new_n204_), .ZN(new_n944_));
  OAI21_X1  g743(.A(G204gat), .B1(new_n934_), .B2(new_n567_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n942_), .B1(new_n944_), .B2(new_n945_), .ZN(G1353gat));
  AOI211_X1 g745(.A(KEYINPUT63), .B(G211gat), .C1(new_n936_), .C2(new_n616_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(KEYINPUT63), .B(G211gat), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n934_), .A2(new_n627_), .A3(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1354gat));
  OR3_X1    g749(.A1(new_n934_), .A2(G218gat), .A3(new_n600_), .ZN(new_n951_));
  OAI21_X1  g750(.A(G218gat), .B1(new_n934_), .B2(new_n899_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1355gat));
endmodule


