//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT77), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n204_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT23), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n210_), .B1(new_n217_), .B2(new_n205_), .ZN(new_n218_));
  OAI22_X1  g017(.A1(new_n216_), .A2(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT79), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G176gat), .ZN(new_n225_));
  INV_X1    g024(.A(G169gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT22), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G169gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n223_), .A2(new_n225_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT80), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT79), .B(G176gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n221_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n219_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G183gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT74), .B1(new_n238_), .B2(KEYINPUT25), .ZN(new_n239_));
  INV_X1    g038(.A(G190gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT26), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G190gat), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n239_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT74), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n238_), .A2(KEYINPUT25), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(G183gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n245_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT24), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n226_), .A3(new_n222_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n244_), .A2(new_n249_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n207_), .A2(new_n209_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n204_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n214_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n206_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n254_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n265_), .A2(KEYINPUT76), .A3(new_n252_), .A4(new_n253_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n255_), .A2(new_n261_), .A3(new_n264_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n237_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G197gat), .B(G204gat), .Z(new_n269_));
  INV_X1    g068(.A(KEYINPUT86), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(KEYINPUT21), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n269_), .A2(KEYINPUT21), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n269_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n203_), .B1(new_n268_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT19), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n216_), .A2(new_n218_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n250_), .A2(KEYINPUT89), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT89), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT24), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n288_), .A2(new_n220_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n254_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT25), .B(G183gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n257_), .A2(new_n260_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n230_), .A2(new_n220_), .ZN(new_n297_));
  OAI22_X1  g096(.A1(new_n284_), .A2(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n280_), .B(new_n283_), .C1(new_n279_), .C2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n203_), .B1(new_n298_), .B2(new_n279_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n237_), .A2(new_n267_), .A3(new_n278_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT90), .B1(new_n302_), .B2(new_n282_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT90), .ZN(new_n304_));
  AOI211_X1 g103(.A(new_n304_), .B(new_n283_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n299_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G8gat), .B(G36gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT92), .ZN(new_n308_));
  XOR2_X1   g107(.A(G64gat), .B(G92gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT93), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n312_), .B(new_n299_), .C1(new_n303_), .C2(new_n305_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n306_), .A2(KEYINPUT93), .A3(new_n313_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321_));
  INV_X1    g120(.A(G141gat), .ZN(new_n322_));
  INV_X1    g121(.A(G148gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(KEYINPUT1), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(G155gat), .A3(G162gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(new_n331_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G141gat), .B(G148gat), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G134gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G127gat), .ZN(new_n343_));
  INV_X1    g142(.A(G127gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G134gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G120gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G113gat), .ZN(new_n348_));
  INV_X1    g147(.A(G113gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G120gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n343_), .A2(new_n345_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n352_), .A2(KEYINPUT85), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT85), .B1(new_n352_), .B2(new_n353_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n341_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n330_), .A2(new_n333_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n353_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n363_));
  NOR2_X1   g162(.A1(new_n356_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n356_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT95), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n356_), .A2(KEYINPUT95), .A3(KEYINPUT4), .A4(new_n359_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n364_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n362_), .B1(new_n369_), .B2(new_n361_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G1gat), .B(G29gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(new_n362_), .C1(new_n369_), .C2(new_n361_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(KEYINPUT100), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT100), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n380_), .A3(new_n375_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n268_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n237_), .A2(new_n267_), .A3(KEYINPUT30), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT31), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT31), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n383_), .A2(new_n384_), .A3(new_n388_), .A4(new_n385_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n355_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n352_), .A2(KEYINPUT85), .A3(new_n353_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n383_), .A2(new_n385_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT84), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT82), .B(KEYINPUT83), .Z(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n398_), .B(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n393_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n384_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n393_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n402_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n390_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n395_), .A2(new_n393_), .A3(new_n402_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n405_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n387_), .A4(new_n389_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n379_), .A2(new_n381_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n302_), .A2(new_n282_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n279_), .B1(new_n298_), .B2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n414_), .B2(new_n298_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n280_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n413_), .B1(new_n417_), .B2(new_n282_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n316_), .B(KEYINPUT27), .C1(new_n418_), .C2(new_n312_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n278_), .B1(KEYINPUT29), .B2(new_n341_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G228gat), .A2(G233gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(KEYINPUT87), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n421_), .B(KEYINPUT87), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n422_), .B(new_n424_), .C1(new_n420_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT88), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n341_), .A2(KEYINPUT29), .ZN(new_n429_));
  XOR2_X1   g228(.A(G22gat), .B(G50gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT28), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n429_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n422_), .B1(new_n420_), .B2(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n423_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n427_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n433_), .A2(new_n436_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n320_), .A2(new_n412_), .A3(new_n419_), .A4(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT101), .ZN(new_n441_));
  INV_X1    g240(.A(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n379_), .A2(new_n381_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n320_), .A2(new_n419_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n312_), .A2(KEYINPUT32), .ZN(new_n447_));
  MUX2_X1   g246(.A(new_n418_), .B(new_n306_), .S(new_n447_), .Z(new_n448_));
  AND3_X1   g247(.A1(new_n448_), .A2(new_n381_), .A3(new_n379_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT94), .B1(new_n317_), .B2(new_n319_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n370_), .A2(KEYINPUT33), .A3(new_n375_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n369_), .A2(new_n361_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n452_), .B(new_n377_), .C1(new_n361_), .C2(new_n360_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT98), .B1(new_n376_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT98), .ZN(new_n457_));
  AOI211_X1 g256(.A(new_n457_), .B(KEYINPUT33), .C1(new_n370_), .C2(new_n375_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n454_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n450_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n317_), .A2(KEYINPUT94), .A3(new_n319_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n449_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n446_), .B1(new_n462_), .B2(new_n442_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n408_), .A2(new_n411_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n441_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT10), .B(G99gat), .Z(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G85gat), .B(G92gat), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT9), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G85gat), .ZN(new_n477_));
  INV_X1    g276(.A(G92gat), .ZN(new_n478_));
  OR3_X1    g277(.A1(new_n477_), .A2(new_n478_), .A3(KEYINPUT9), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n469_), .A2(new_n471_), .A3(new_n476_), .A4(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G29gat), .B(G36gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT67), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n483_));
  INV_X1    g282(.A(G29gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(G36gat), .ZN(new_n485_));
  INV_X1    g284(.A(G36gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(G29gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n483_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n482_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n474_), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT64), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT64), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n473_), .A2(new_n475_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n493_), .B1(new_n503_), .B2(new_n470_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n470_), .A2(new_n493_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n476_), .B2(new_n502_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n480_), .B(new_n492_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT34), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n507_), .A2(KEYINPUT69), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT69), .B1(new_n507_), .B2(new_n512_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n480_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT66), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n518_), .B(new_n480_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n492_), .A2(KEYINPUT15), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT68), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n517_), .A2(KEYINPUT68), .A3(new_n519_), .A4(new_n523_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n515_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n510_), .A2(new_n511_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G190gat), .B(G218gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT36), .ZN(new_n534_));
  INV_X1    g333(.A(new_n529_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n507_), .A2(new_n535_), .A3(new_n512_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n524_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n524_), .A2(new_n536_), .A3(KEYINPUT70), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n530_), .A2(new_n534_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n533_), .B(KEYINPUT36), .Z(new_n544_));
  AND3_X1   g343(.A1(new_n530_), .A2(KEYINPUT71), .A3(new_n541_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT71), .B1(new_n530_), .B2(new_n541_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(KEYINPUT72), .B(new_n544_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n543_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT73), .B(G15gat), .ZN(new_n552_));
  INV_X1    g351(.A(G22gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n558_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n564_));
  XOR2_X1   g363(.A(G71gat), .B(G78gat), .Z(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n564_), .A2(new_n565_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n562_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G155gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n573_), .A2(new_n574_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(KEYINPUT17), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n573_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT65), .B1(new_n516_), .B2(new_n569_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n516_), .B2(new_n569_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n516_), .A2(KEYINPUT65), .A3(new_n569_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(G230gat), .A3(G233gat), .A4(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT12), .B1(new_n516_), .B2(new_n569_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n516_), .A2(new_n569_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n569_), .A2(KEYINPUT12), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n517_), .A2(new_n519_), .A3(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n590_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT5), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G176gat), .B(G204gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n586_), .A2(new_n594_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT13), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(KEYINPUT13), .A3(new_n602_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n492_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n562_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n560_), .A2(new_n492_), .A3(new_n561_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n562_), .A2(new_n523_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n611_), .A2(new_n608_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G169gat), .B(G197gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n614_), .A2(new_n613_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n612_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n607_), .A2(new_n623_), .ZN(new_n624_));
  NOR4_X1   g423(.A1(new_n466_), .A2(new_n551_), .A3(new_n582_), .A4(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n443_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n202_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT102), .ZN(new_n628_));
  INV_X1    g427(.A(new_n623_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n582_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n543_), .A2(KEYINPUT37), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n530_), .A2(new_n541_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n544_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n636_), .B2(new_n542_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n607_), .B(new_n630_), .C1(new_n633_), .C2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n466_), .A2(new_n629_), .A3(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n202_), .A3(new_n626_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT38), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n628_), .A2(new_n641_), .ZN(G1324gat));
  AOI21_X1  g441(.A(new_n555_), .B1(new_n625_), .B2(new_n445_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT39), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n639_), .A2(new_n555_), .A3(new_n445_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(G1325gat));
  INV_X1    g447(.A(G15gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n625_), .B2(new_n464_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT41), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n639_), .A2(new_n649_), .A3(new_n464_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1326gat));
  AOI21_X1  g452(.A(new_n553_), .B1(new_n625_), .B2(new_n442_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT42), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n639_), .A2(new_n553_), .A3(new_n442_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n466_), .A2(new_n629_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n551_), .A2(new_n582_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n607_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n626_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT71), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n635_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n530_), .A2(KEYINPUT71), .A3(new_n541_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT72), .B1(new_n669_), .B2(new_n544_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n550_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n631_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n637_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n317_), .A2(new_n319_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT94), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n451_), .A2(new_n453_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n376_), .A2(new_n455_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n457_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n376_), .A2(KEYINPUT98), .A3(new_n455_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n677_), .A2(new_n682_), .A3(new_n461_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n626_), .A2(new_n448_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n442_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n444_), .A2(new_n445_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n465_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n440_), .B(KEYINPUT101), .Z(new_n688_));
  AOI21_X1  g487(.A(new_n674_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n665_), .B1(new_n689_), .B2(KEYINPUT103), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n691_), .B(KEYINPUT43), .C1(new_n466_), .C2(new_n674_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n630_), .A2(new_n624_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT44), .B1(new_n693_), .B2(new_n694_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n443_), .A2(new_n484_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n664_), .B1(new_n697_), .B2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n445_), .B(KEYINPUT104), .Z(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n662_), .A2(KEYINPUT105), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT105), .B1(new_n662_), .B2(new_n703_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(KEYINPUT45), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT45), .B1(new_n704_), .B2(new_n705_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n486_), .B1(new_n697_), .B2(new_n445_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT106), .B(new_n700_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n700_), .A2(KEYINPUT106), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n706_), .A2(new_n707_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n697_), .A2(new_n445_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n711_), .B(new_n712_), .C1(new_n713_), .C2(new_n486_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(G1329gat));
  AOI21_X1  g514(.A(G43gat), .B1(new_n663_), .B2(new_n464_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n464_), .A2(G43gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n697_), .B2(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g518(.A(G50gat), .B1(new_n663_), .B2(new_n442_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n442_), .A2(G50gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n697_), .B2(new_n721_), .ZN(G1331gat));
  NAND3_X1  g521(.A1(new_n630_), .A2(new_n629_), .A3(new_n660_), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n466_), .A2(new_n551_), .A3(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT107), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(G57gat), .A3(new_n626_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT108), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT108), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n466_), .A2(new_n623_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n582_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n660_), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n626_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n727_), .A2(new_n728_), .A3(new_n733_), .ZN(G1332gat));
  INV_X1    g533(.A(G64gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n701_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n725_), .B2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT48), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n732_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n725_), .B2(new_n464_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT49), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n464_), .A2(new_n741_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT109), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n731_), .B2(new_n745_), .ZN(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n725_), .B2(new_n442_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT50), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n732_), .A2(new_n747_), .A3(new_n442_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1335gat));
  NOR3_X1   g550(.A1(new_n630_), .A2(new_n623_), .A3(new_n607_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT110), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT110), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n443_), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n466_), .A2(new_n623_), .A3(new_n607_), .A4(new_n659_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n477_), .A3(new_n626_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1336gat));
  OAI21_X1  g560(.A(G92gat), .B1(new_n757_), .B2(new_n701_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n478_), .A3(new_n445_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n467_), .A3(new_n464_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(KEYINPUT111), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n464_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G99gat), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n766_), .A2(KEYINPUT111), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n759_), .A2(new_n468_), .A3(new_n442_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n439_), .B(new_n753_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n468_), .B1(new_n775_), .B2(KEYINPUT112), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT112), .B1(new_n754_), .B2(new_n442_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n774_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n693_), .A2(KEYINPUT112), .A3(new_n442_), .A4(new_n752_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G106gat), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(new_n777_), .A3(new_n773_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n772_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n772_), .C1(new_n779_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT54), .B1(new_n638_), .B2(new_n623_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n730_), .A2(new_n790_), .A3(new_n629_), .A4(new_n607_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n590_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n594_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n589_), .A2(new_n593_), .A3(KEYINPUT55), .A4(new_n590_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n599_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n800_), .B(new_n601_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n623_), .A2(new_n602_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n610_), .A2(new_n611_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n618_), .B1(new_n804_), .B2(new_n608_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n611_), .A2(new_n613_), .A3(G229gat), .A4(G233gat), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n615_), .A2(new_n618_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n802_), .A2(new_n803_), .B1(new_n603_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n793_), .B1(new_n551_), .B2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n807_), .A2(new_n602_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n810_), .B(KEYINPUT58), .C1(new_n799_), .C2(new_n801_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n809_), .B1(new_n674_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n542_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n803_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n603_), .A2(new_n807_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(KEYINPUT57), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n817_), .A2(KEYINPUT114), .A3(new_n820_), .A4(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n816_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n792_), .B1(new_n825_), .B2(new_n630_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n445_), .A2(new_n442_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n626_), .A3(new_n464_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n788_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n815_), .A2(new_n633_), .A3(new_n637_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n817_), .B2(new_n820_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT115), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n823_), .A2(new_n824_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n809_), .B(new_n835_), .C1(new_n674_), .C2(new_n815_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n582_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(KEYINPUT116), .A3(new_n582_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n792_), .A3(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n828_), .A2(KEYINPUT59), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n830_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n349_), .B1(new_n844_), .B2(new_n623_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n792_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n831_), .A2(new_n832_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n630_), .B1(new_n834_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n828_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n349_), .A3(new_n623_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n845_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n629_), .B(new_n830_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n854_), .B(new_n851_), .C1(new_n855_), .C2(new_n349_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1340gat));
  OAI21_X1  g656(.A(new_n347_), .B1(new_n607_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n850_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n347_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT118), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n844_), .A2(new_n660_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n347_), .ZN(G1341gat));
  NAND3_X1  g661(.A1(new_n850_), .A2(new_n344_), .A3(new_n630_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n844_), .A2(new_n630_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n344_), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n850_), .B2(new_n551_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n674_), .A2(new_n342_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT119), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n844_), .B2(new_n868_), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n849_), .A2(new_n464_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n736_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n629_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n322_), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n607_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n323_), .ZN(G1345gat));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n872_), .B2(new_n582_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n870_), .A2(KEYINPUT120), .A3(new_n630_), .A4(new_n871_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n872_), .A2(new_n884_), .A3(new_n674_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n872_), .B2(new_n817_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n887_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1347gat));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n736_), .A2(new_n412_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n439_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n623_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n846_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n841_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n891_), .B1(new_n898_), .B2(new_n226_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n837_), .A2(KEYINPUT116), .A3(new_n582_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT116), .B1(new_n837_), .B2(new_n582_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n900_), .A2(new_n901_), .A3(new_n846_), .ZN(new_n902_));
  OAI211_X1 g701(.A(KEYINPUT62), .B(G169gat), .C1(new_n902_), .C2(new_n896_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n898_), .A2(new_n233_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n899_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT122), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n899_), .A2(new_n903_), .A3(new_n907_), .A4(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1348gat));
  INV_X1    g708(.A(new_n232_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n894_), .B1(new_n897_), .B2(new_n841_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n660_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT123), .B1(new_n849_), .B2(new_n442_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n826_), .A2(new_n914_), .A3(new_n439_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n607_), .A2(new_n222_), .ZN(new_n916_));
  AND4_X1   g715(.A1(new_n893_), .A2(new_n913_), .A3(new_n915_), .A4(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n912_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT124), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n912_), .B2(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1349gat));
  INV_X1    g721(.A(new_n911_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n923_), .A2(new_n292_), .A3(new_n582_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n913_), .A2(new_n630_), .A3(new_n893_), .A4(new_n915_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n238_), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n923_), .B2(new_n674_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n911_), .A2(new_n551_), .A3(new_n293_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1351gat));
  NOR2_X1   g728(.A1(new_n701_), .A2(new_n444_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n465_), .B(new_n930_), .C1(new_n846_), .C2(new_n848_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n623_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g733(.A(G204gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n660_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n932_), .A2(KEYINPUT125), .A3(new_n660_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT126), .B1(new_n936_), .B2(G204gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n940_), .B2(new_n938_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1353gat));
  NOR2_X1   g743(.A1(new_n931_), .A2(new_n582_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT63), .B(G211gat), .Z(new_n946_));
  AOI21_X1  g745(.A(KEYINPUT127), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  MUX2_X1   g747(.A(new_n948_), .B(new_n946_), .S(new_n945_), .Z(new_n949_));
  AOI21_X1  g748(.A(new_n947_), .B1(new_n949_), .B2(KEYINPUT127), .ZN(G1354gat));
  OAI21_X1  g749(.A(G218gat), .B1(new_n931_), .B2(new_n674_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n817_), .A2(G218gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n931_), .B2(new_n952_), .ZN(G1355gat));
endmodule


