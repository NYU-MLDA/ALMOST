//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .A4(KEYINPUT65), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n218_), .A2(new_n220_), .B1(new_n221_), .B2(KEYINPUT8), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n221_), .A2(KEYINPUT8), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n216_), .B(new_n222_), .C1(new_n221_), .C2(KEYINPUT8), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n217_), .B1(new_n227_), .B2(new_n219_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT64), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n231_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n219_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n205_), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n213_), .A3(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n225_), .A2(new_n226_), .A3(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G29gat), .B(G36gat), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n240_), .A2(KEYINPUT70), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(KEYINPUT70), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n239_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n238_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n234_), .A2(KEYINPUT67), .A3(new_n213_), .A4(new_n237_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n225_), .A2(new_n226_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT15), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n246_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT15), .A3(new_n244_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT34), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT35), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n248_), .A2(new_n257_), .A3(new_n258_), .A4(new_n263_), .ZN(new_n264_));
  AOI211_X1 g063(.A(new_n262_), .B(new_n261_), .C1(new_n257_), .C2(KEYINPUT71), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n262_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n248_), .A2(new_n257_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n264_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT73), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G190gat), .B(G218gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G134gat), .B(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT36), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT72), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n268_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n273_), .A2(KEYINPUT36), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n270_), .A2(new_n277_), .B1(new_n278_), .B2(new_n268_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G43gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(G15gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT23), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(G183gat), .A3(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT24), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n295_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT26), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n301_));
  INV_X1    g100(.A(G183gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(KEYINPUT25), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(KEYINPUT25), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT25), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n300_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n288_), .B2(new_n286_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(new_n288_), .B2(new_n286_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT82), .B(G176gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n295_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n297_), .A2(new_n306_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT30), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT83), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n315_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n285_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n317_), .A2(new_n285_), .ZN(new_n319_));
  INV_X1    g118(.A(G134gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G127gat), .ZN(new_n321_));
  INV_X1    g120(.A(G127gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G134gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT84), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n323_), .A3(KEYINPUT84), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n321_), .A2(new_n323_), .A3(KEYINPUT84), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(new_n324_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OR3_X1    g134(.A1(new_n318_), .A2(new_n319_), .A3(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT86), .Z(new_n339_));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342_));
  AND2_X1   g141(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n343_), .A2(new_n344_), .A3(G197gat), .ZN(new_n345_));
  INV_X1    g144(.A(G197gat), .ZN(new_n346_));
  INV_X1    g145(.A(G204gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT21), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n342_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(G197gat), .B1(new_n343_), .B2(new_n344_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT21), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT93), .B1(new_n349_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT21), .ZN(new_n355_));
  OR2_X1    g154(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n346_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n355_), .B1(new_n358_), .B2(new_n351_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  INV_X1    g159(.A(G218gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G211gat), .ZN(new_n362_));
  INV_X1    g161(.A(G211gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G218gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n346_), .A3(new_n357_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n355_), .B1(G197gat), .B2(G204gat), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n359_), .A2(new_n360_), .A3(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n350_), .A2(new_n365_), .A3(KEYINPUT21), .A4(new_n352_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT94), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n342_), .A2(new_n355_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n352_), .A4(new_n350_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n354_), .A2(new_n369_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT89), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n379_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT88), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n387_), .A2(KEYINPUT88), .A3(new_n388_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n381_), .B(new_n386_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n391_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n395_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT1), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n394_), .A2(new_n405_), .A3(new_n395_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n406_), .A3(new_n398_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n382_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n387_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n376_), .B1(new_n401_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n341_), .B1(new_n375_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n371_), .A2(new_n374_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n349_), .A2(new_n353_), .A3(KEYINPUT93), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n360_), .B1(new_n359_), .B2(new_n368_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n384_), .A2(new_n385_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n389_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n387_), .A2(KEYINPUT88), .A3(new_n388_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n399_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n409_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n397_), .B1(new_n396_), .B2(KEYINPUT1), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n406_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT29), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n416_), .A2(new_n340_), .A3(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n412_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n412_), .A2(new_n427_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT96), .B1(new_n433_), .B2(new_n428_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT96), .ZN(new_n435_));
  AOI211_X1 g234(.A(new_n435_), .B(new_n429_), .C1(new_n412_), .C2(new_n427_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n438_));
  AOI22_X1  g237(.A1(new_n391_), .A2(new_n400_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT90), .A3(new_n376_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT90), .B1(new_n439_), .B2(new_n376_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n438_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G22gat), .B(G50gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n446_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n447_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n432_), .A2(new_n437_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n433_), .A2(new_n428_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n448_), .A3(new_n453_), .A4(new_n430_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(G85gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT0), .B(G57gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT101), .B(new_n332_), .C1(new_n422_), .C2(new_n425_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n401_), .A2(new_n410_), .A3(new_n328_), .A4(new_n331_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT4), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n401_), .A2(new_n410_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(KEYINPUT101), .A3(new_n468_), .A4(new_n332_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n463_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n463_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n401_), .A2(new_n410_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n473_), .B2(new_n465_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n462_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n470_), .A2(new_n462_), .A3(new_n474_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT18), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G64gat), .B(G92gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n483_), .A2(KEYINPUT32), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n309_), .A2(new_n312_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT98), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n299_), .A2(G190gat), .ZN(new_n487_));
  INV_X1    g286(.A(G190gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(KEYINPUT26), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(KEYINPUT26), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n299_), .A2(G190gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT98), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT25), .B(G183gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n296_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT99), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n294_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n290_), .A2(KEYINPUT99), .A3(new_n293_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n485_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT20), .B1(new_n375_), .B2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n313_), .B(new_n413_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G226gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n502_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n375_), .B2(new_n501_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n313_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n416_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n507_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n484_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n508_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n513_), .A3(new_n507_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n515_), .B1(new_n518_), .B2(new_n484_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n478_), .A2(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n516_), .A2(new_n483_), .A3(new_n517_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n483_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT100), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n475_), .A2(KEYINPUT33), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n525_), .B(new_n462_), .C1(new_n470_), .C2(new_n474_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n465_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(new_n472_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n462_), .B1(new_n529_), .B2(new_n471_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n466_), .A2(KEYINPUT102), .A3(new_n463_), .A4(new_n469_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n466_), .A2(new_n463_), .A3(new_n469_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT102), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n511_), .A2(new_n513_), .A3(new_n507_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT98), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT98), .B1(new_n491_), .B2(new_n492_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n495_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n296_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n499_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT99), .B1(new_n290_), .B2(new_n293_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n540_), .B(new_n541_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n485_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n510_), .B1(new_n416_), .B2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n507_), .B1(new_n547_), .B2(new_n503_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n482_), .B1(new_n537_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT100), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n516_), .A2(new_n483_), .A3(new_n517_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n523_), .A2(new_n527_), .A3(new_n536_), .A4(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT103), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n520_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n524_), .A2(new_n526_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n556_), .A2(KEYINPUT103), .A3(new_n523_), .A4(new_n552_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n457_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n478_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT27), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n551_), .A2(KEYINPUT104), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT104), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n516_), .A2(new_n562_), .A3(new_n517_), .A4(new_n483_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n482_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n560_), .B1(KEYINPUT27), .B2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n559_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n339_), .B1(new_n558_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n566_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n338_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(new_n478_), .A3(new_n456_), .A4(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n279_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT106), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(new_n573_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT11), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n580_));
  INV_X1    g379(.A(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n579_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT74), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G15gat), .B(G22gat), .ZN(new_n588_));
  INV_X1    g387(.A(G8gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G1gat), .B(G8gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n587_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT17), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n599_), .A2(new_n600_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n595_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT75), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n225_), .A2(new_n584_), .A3(new_n226_), .A4(new_n238_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT12), .ZN(new_n608_));
  INV_X1    g407(.A(new_n584_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n239_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT12), .B(new_n579_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n252_), .A2(KEYINPUT68), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT68), .B1(new_n252_), .B2(new_n614_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n611_), .B(new_n612_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n610_), .A2(new_n607_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n612_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT5), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n621_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT13), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n627_), .B1(KEYINPUT69), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n255_), .A2(new_n244_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT76), .B1(new_n633_), .B2(new_n593_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(KEYINPUT76), .A3(new_n593_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT77), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G229gat), .A2(G233gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n254_), .A2(new_n256_), .A3(new_n594_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .A4(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n636_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n640_), .B(new_n639_), .C1(new_n642_), .C2(new_n634_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT77), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n247_), .A2(new_n594_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n639_), .B1(new_n637_), .B2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT79), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G169gat), .B(G197gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(KEYINPUT78), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n647_), .A2(new_n653_), .ZN(new_n654_));
  OAI221_X1 g453(.A(new_n641_), .B1(KEYINPUT78), .B2(new_n652_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n632_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n606_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n576_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n478_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n202_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n553_), .A2(new_n554_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n520_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n557_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n567_), .B1(new_n666_), .B2(new_n456_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n338_), .B(KEYINPUT86), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n571_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n657_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT105), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n270_), .A2(new_n277_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n268_), .A2(new_n278_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT37), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n673_), .B(KEYINPUT37), .C1(new_n268_), .C2(new_n275_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n605_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n632_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n671_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n202_), .A3(new_n661_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n662_), .B1(new_n663_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(new_n663_), .B2(new_n682_), .ZN(G1324gat));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n589_), .A3(new_n566_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n566_), .B(new_n659_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT39), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G8gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G8gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1325gat));
  NAND3_X1  g491(.A1(new_n681_), .A2(new_n283_), .A3(new_n668_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n660_), .A2(new_n668_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n694_), .B2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1326gat));
  INV_X1    g496(.A(G22gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n681_), .A2(new_n698_), .A3(new_n457_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n660_), .A2(new_n457_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(G22gat), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT42), .B(new_n698_), .C1(new_n660_), .C2(new_n457_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1327gat));
  NOR2_X1   g503(.A1(new_n658_), .A2(new_n605_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT107), .B(new_n675_), .C1(new_n279_), .C2(KEYINPUT37), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n706_), .B1(new_n669_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n677_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n706_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT44), .B(new_n705_), .C1(new_n712_), .C2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n669_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n710_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n706_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT44), .B1(new_n721_), .B2(new_n705_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n717_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724_), .B2(new_n478_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n279_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n605_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT108), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n679_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n671_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G29gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n661_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n725_), .A2(new_n732_), .ZN(G1328gat));
  NOR2_X1   g532(.A1(new_n569_), .A2(G36gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n671_), .A2(new_n729_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT45), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n671_), .A2(new_n737_), .A3(new_n729_), .A4(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n723_), .B2(new_n566_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n705_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n745_), .A2(new_n741_), .A3(new_n566_), .A4(new_n716_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G36gat), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n739_), .B(new_n740_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n566_), .A3(new_n716_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT109), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(G36gat), .A3(new_n746_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n740_), .B1(new_n752_), .B2(new_n739_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n749_), .A2(new_n753_), .ZN(G1329gat));
  NAND3_X1  g553(.A1(new_n723_), .A2(G43gat), .A3(new_n570_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n671_), .A2(new_n668_), .A3(new_n729_), .ZN(new_n756_));
  INV_X1    g555(.A(G43gat), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(KEYINPUT111), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT111), .B1(new_n756_), .B2(new_n757_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT47), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n755_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1330gat));
  AOI21_X1  g563(.A(G50gat), .B1(new_n730_), .B2(new_n457_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n457_), .A2(G50gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n723_), .B2(new_n766_), .ZN(G1331gat));
  NAND2_X1  g566(.A1(new_n679_), .A2(new_n656_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n606_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n576_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n661_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G57gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n657_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n678_), .A2(new_n632_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(G57gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n661_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n776_), .B2(new_n778_), .ZN(G1332gat));
  OR3_X1    g578(.A1(new_n776_), .A2(G64gat), .A3(new_n569_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G64gat), .B1(new_n770_), .B2(new_n569_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n782_), .B2(new_n783_), .ZN(G1333gat));
  OR3_X1    g583(.A1(new_n776_), .A2(G71gat), .A3(new_n339_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n771_), .A2(new_n668_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(G71gat), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G71gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1334gat));
  OR3_X1    g589(.A1(new_n776_), .A2(G78gat), .A3(new_n456_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n457_), .B(new_n769_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(G78gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G78gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT113), .ZN(G1335gat));
  NAND2_X1  g596(.A1(new_n669_), .A2(new_n656_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n728_), .A2(new_n798_), .A3(new_n632_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n219_), .A3(new_n661_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n768_), .A2(new_n605_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n721_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n661_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n804_), .B2(new_n219_), .ZN(G1336gat));
  AOI21_X1  g604(.A(new_n217_), .B1(new_n802_), .B2(new_n566_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n799_), .A2(new_n217_), .A3(new_n566_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT114), .ZN(G1337gat));
  NAND4_X1  g608(.A1(new_n799_), .A2(new_n570_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n802_), .A2(new_n668_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n812_), .B2(new_n204_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g613(.A1(new_n799_), .A2(new_n205_), .A3(new_n457_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n721_), .A2(new_n457_), .A3(new_n801_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(G106gat), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(G106gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n815_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n569_), .A2(new_n456_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n570_), .A2(new_n661_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n647_), .A2(new_n652_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  INV_X1    g626(.A(new_n639_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n640_), .B(new_n828_), .C1(new_n642_), .C2(new_n634_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n651_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n637_), .B2(new_n645_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n645_), .B1(new_n642_), .B2(new_n634_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n639_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(KEYINPUT118), .A3(new_n651_), .A4(new_n829_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n826_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n627_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n617_), .A2(new_n620_), .A3(new_n626_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n654_), .A2(new_n655_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n252_), .A2(new_n614_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT68), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n252_), .A2(KEYINPUT68), .A3(new_n614_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n612_), .B1(new_n846_), .B2(new_n611_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n617_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n611_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n850_), .A2(new_n848_), .A3(new_n619_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n841_), .B(new_n626_), .C1(new_n849_), .C2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n840_), .B1(new_n853_), .B2(KEYINPUT116), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n848_), .B1(new_n850_), .B2(new_n619_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n617_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n625_), .B1(new_n857_), .B2(new_n851_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n841_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT56), .B(new_n625_), .C1(new_n857_), .C2(new_n851_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n854_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n838_), .B1(new_n863_), .B2(KEYINPUT117), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n854_), .A2(new_n862_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n279_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n826_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n826_), .A2(new_n836_), .A3(new_n870_), .A4(new_n839_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n859_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n872_), .B(KEYINPUT58), .C1(new_n853_), .C2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n853_), .B2(new_n873_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n677_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n867_), .A2(KEYINPUT57), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879_));
  INV_X1    g678(.A(new_n866_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n865_), .B1(new_n854_), .B2(new_n862_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n880_), .A2(new_n881_), .A3(new_n838_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n882_), .B2(new_n279_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n605_), .B1(new_n878_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n680_), .A2(new_n656_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n885_), .A2(KEYINPUT54), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(KEYINPUT54), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n822_), .B(new_n825_), .C1(new_n884_), .C2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT119), .B1(new_n867_), .B2(KEYINPUT57), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n891_), .B(new_n879_), .C1(new_n882_), .C2(new_n279_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n878_), .A2(new_n890_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n888_), .B1(new_n893_), .B2(new_n606_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n825_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n657_), .B(new_n889_), .C1(new_n896_), .C2(new_n822_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G113gat), .ZN(new_n898_));
  INV_X1    g697(.A(G113gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n899_), .A3(new_n657_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1340gat));
  OAI211_X1 g700(.A(new_n679_), .B(new_n889_), .C1(new_n896_), .C2(new_n822_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G120gat), .ZN(new_n903_));
  INV_X1    g702(.A(G120gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n632_), .B2(KEYINPUT60), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n896_), .B(new_n905_), .C1(KEYINPUT60), .C2(new_n904_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(G1341gat));
  OAI211_X1 g706(.A(new_n605_), .B(new_n889_), .C1(new_n896_), .C2(new_n822_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G127gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n896_), .A2(new_n322_), .A3(new_n605_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1342gat));
  NAND2_X1  g710(.A1(new_n896_), .A2(new_n279_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n320_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT121), .B(G134gat), .Z(new_n914_));
  NOR2_X1   g713(.A1(new_n677_), .A2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n889_), .B(new_n915_), .C1(new_n896_), .C2(new_n822_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n913_), .A2(new_n916_), .ZN(G1343gat));
  NAND4_X1  g716(.A1(new_n339_), .A2(new_n661_), .A3(new_n457_), .A4(new_n569_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n894_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n657_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n679_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(G148gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1345gat));
  NAND2_X1  g723(.A1(new_n919_), .A2(new_n605_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT61), .B(G155gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1346gat));
  AOI21_X1  g726(.A(G162gat), .B1(new_n919_), .B2(new_n279_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n711_), .A2(G162gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n919_), .B2(new_n929_), .ZN(G1347gat));
  NOR3_X1   g729(.A1(new_n339_), .A2(new_n661_), .A3(new_n569_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n456_), .B(new_n931_), .C1(new_n884_), .C2(new_n888_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G169gat), .B1(new_n932_), .B2(new_n656_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n867_), .A2(KEYINPUT57), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n877_), .A2(new_n874_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n867_), .A2(KEYINPUT57), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n606_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n886_), .A2(new_n887_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n457_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n942_), .A2(new_n311_), .A3(new_n657_), .A4(new_n931_), .ZN(new_n943_));
  OAI211_X1 g742(.A(KEYINPUT62), .B(G169gat), .C1(new_n932_), .C2(new_n656_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n935_), .A2(new_n943_), .A3(new_n944_), .ZN(G1348gat));
  NAND3_X1  g744(.A1(new_n931_), .A2(G176gat), .A3(new_n679_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n894_), .A2(new_n457_), .A3(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n310_), .B1(new_n932_), .B2(new_n632_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(KEYINPUT123), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n950_), .B(new_n310_), .C1(new_n932_), .C2(new_n632_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n947_), .B1(new_n949_), .B2(new_n951_), .ZN(G1349gat));
  NAND2_X1  g751(.A1(new_n931_), .A2(new_n605_), .ZN(new_n953_));
  OR3_X1    g752(.A1(new_n894_), .A2(new_n457_), .A3(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n495_), .ZN(new_n955_));
  AOI22_X1  g754(.A1(new_n954_), .A2(new_n302_), .B1(new_n942_), .B2(new_n955_), .ZN(G1350gat));
  NAND4_X1  g755(.A1(new_n942_), .A2(new_n494_), .A3(new_n279_), .A4(new_n931_), .ZN(new_n957_));
  OAI21_X1  g756(.A(G190gat), .B1(new_n932_), .B2(new_n677_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n957_), .A2(new_n958_), .A3(KEYINPUT124), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1351gat));
  NAND4_X1  g762(.A1(new_n339_), .A2(new_n478_), .A3(new_n457_), .A4(new_n566_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n893_), .A2(new_n606_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n964_), .B1(new_n965_), .B2(new_n941_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n657_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n356_), .A2(new_n357_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  AND4_X1   g770(.A1(new_n969_), .A2(new_n966_), .A3(new_n971_), .A4(new_n679_), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n894_), .A2(new_n632_), .A3(new_n964_), .ZN(new_n973_));
  OR2_X1    g772(.A1(new_n973_), .A2(new_n347_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n969_), .B1(new_n973_), .B2(new_n971_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n972_), .B1(new_n974_), .B2(new_n975_), .ZN(G1353gat));
  AOI21_X1  g775(.A(new_n606_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n966_), .A2(new_n977_), .ZN(new_n978_));
  OR2_X1    g777(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n979_));
  XNOR2_X1  g778(.A(new_n978_), .B(new_n979_), .ZN(G1354gat));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n361_), .B1(new_n966_), .B2(new_n713_), .ZN(new_n982_));
  NOR4_X1   g781(.A1(new_n894_), .A2(G218gat), .A3(new_n726_), .A4(new_n964_), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n981_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n966_), .A2(new_n361_), .A3(new_n279_), .ZN(new_n985_));
  NOR3_X1   g784(.A1(new_n894_), .A2(new_n677_), .A3(new_n964_), .ZN(new_n986_));
  OAI211_X1 g785(.A(new_n985_), .B(KEYINPUT126), .C1(new_n986_), .C2(new_n361_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n984_), .A2(new_n987_), .ZN(G1355gat));
endmodule


