//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT93), .ZN(new_n204_));
  XOR2_X1   g003(.A(G64gat), .B(G92gat), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n206_), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n207_), .A2(KEYINPUT32), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G226gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT19), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT22), .B(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT23), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  INV_X1    g022(.A(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n217_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(new_n216_), .A3(KEYINPUT80), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(G169gat), .B2(G176gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n229_), .A2(new_n231_), .A3(KEYINPUT24), .A4(new_n213_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n223_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT26), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n238_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT26), .B(G190gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n240_), .B2(KEYINPUT79), .ZN(new_n241_));
  OAI211_X1 g040(.A(KEYINPUT81), .B(new_n232_), .C1(new_n237_), .C2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT24), .B1(new_n229_), .B2(new_n231_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n220_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n221_), .A2(new_n245_), .B1(KEYINPUT23), .B2(new_n218_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G183gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n251_), .A3(new_n235_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n233_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n224_), .A2(KEYINPUT26), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n238_), .A2(G190gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT79), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n238_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT81), .B1(new_n259_), .B2(new_n232_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n227_), .B1(new_n248_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G218gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G211gat), .ZN(new_n266_));
  INV_X1    g065(.A(G211gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G218gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT89), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n264_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(G197gat), .A2(G204gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n273_), .A2(KEYINPUT90), .A3(KEYINPUT21), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n264_), .B(new_n275_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n261_), .A2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n246_), .A2(new_n244_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n217_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n249_), .A2(new_n251_), .A3(new_n254_), .A4(new_n255_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n232_), .A2(new_n283_), .A3(new_n222_), .ZN(new_n284_));
  OAI22_X1  g083(.A1(new_n281_), .A2(new_n282_), .B1(new_n284_), .B2(new_n243_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n212_), .B1(new_n280_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n233_), .A2(new_n252_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n232_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n277_), .A2(new_n278_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n227_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n279_), .B2(new_n285_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n296_), .A2(new_n212_), .A3(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n209_), .B(KEYINPUT97), .C1(new_n289_), .C2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G141gat), .B(G148gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(KEYINPUT1), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n304_), .B2(KEYINPUT1), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT85), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n306_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n301_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G155gat), .B(G162gat), .Z(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  INV_X1    g114(.A(G141gat), .ZN(new_n316_));
  INV_X1    g115(.A(G148gat), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .A4(KEYINPUT86), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n319_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(KEYINPUT3), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n318_), .A2(new_n320_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n311_), .B1(new_n314_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n310_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n310_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n310_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n328_), .B1(new_n310_), .B2(new_n324_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n325_), .A2(new_n336_), .A3(new_n329_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n333_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT0), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n342_), .A2(KEYINPUT0), .ZN(new_n345_));
  OAI21_X1  g144(.A(G57gat), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G1gat), .B(G29gat), .Z(new_n347_));
  INV_X1    g146(.A(KEYINPUT0), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G57gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n343_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n346_), .A2(G85gat), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(G85gat), .B1(new_n346_), .B2(new_n351_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n341_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n352_), .A2(new_n353_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n356_), .B(new_n333_), .C1(new_n337_), .C2(new_n340_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n204_), .B(new_n205_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n296_), .A2(new_n298_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n211_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n211_), .A2(new_n297_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT92), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n286_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT92), .B1(new_n279_), .B2(new_n285_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n280_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n300_), .A2(new_n358_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n296_), .A2(new_n212_), .A3(new_n298_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n295_), .B1(new_n294_), .B2(new_n227_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n372_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n373_), .B2(new_n212_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT97), .B1(new_n374_), .B2(new_n209_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n207_), .A2(new_n208_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n232_), .A2(new_n222_), .A3(new_n283_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n243_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n221_), .A2(new_n245_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n219_), .A3(new_n244_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n225_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n377_), .A2(new_n378_), .B1(new_n381_), .B2(new_n217_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(new_n365_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(new_n367_), .A3(new_n363_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n372_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n212_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n376_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n330_), .A2(new_n331_), .A3(new_n339_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n388_), .A2(new_n354_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n388_), .B2(new_n354_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n338_), .A2(new_n332_), .ZN(new_n392_));
  OAI22_X1  g191(.A1(new_n390_), .A2(new_n391_), .B1(new_n337_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n362_), .A2(new_n368_), .A3(new_n359_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n357_), .B(new_n396_), .ZN(new_n397_));
  OAI22_X1  g196(.A1(new_n370_), .A2(new_n375_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n399_));
  NAND2_X1  g198(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(G228gat), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n310_), .B2(new_n324_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n295_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n312_), .B(KEYINPUT87), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n318_), .A2(new_n322_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n320_), .A2(new_n321_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(G155gat), .B2(G162gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT85), .B1(new_n413_), .B2(new_n302_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n308_), .B1(new_n414_), .B2(new_n303_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n411_), .A2(new_n311_), .B1(new_n415_), .B2(new_n301_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n279_), .B(new_n403_), .C1(new_n416_), .C2(new_n405_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n407_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n407_), .B2(new_n417_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n399_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n295_), .A2(new_n406_), .A3(new_n404_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n325_), .A2(KEYINPUT29), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n403_), .B1(new_n424_), .B2(new_n279_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n407_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(KEYINPUT91), .A3(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G22gat), .B(G50gat), .Z(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT28), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n325_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n429_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n422_), .A2(new_n428_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n436_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n439_), .A2(KEYINPUT91), .A3(new_n427_), .A4(new_n426_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n398_), .A2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n438_), .A2(new_n440_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n358_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n385_), .A2(new_n376_), .A3(new_n386_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n359_), .B1(new_n362_), .B2(new_n368_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n376_), .B1(new_n289_), .B2(new_n299_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n394_), .A3(KEYINPUT27), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n443_), .A2(new_n444_), .A3(new_n448_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n442_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(G15gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(G71gat), .B(G99gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(G43gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n294_), .A2(new_n227_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n294_), .B2(new_n227_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT31), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n261_), .A2(new_n459_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n458_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n294_), .A2(new_n227_), .A3(new_n460_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n463_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n464_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n329_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n461_), .A2(new_n462_), .A3(new_n458_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n466_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT31), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n463_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n328_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n452_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT98), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n328_), .A3(new_n475_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n329_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n441_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n448_), .A2(new_n444_), .A3(new_n450_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n480_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n449_), .A2(KEYINPUT27), .A3(new_n394_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT27), .B1(new_n387_), .B2(new_n394_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n358_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(KEYINPUT98), .A3(new_n477_), .A4(new_n441_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n479_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G29gat), .B(G36gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500_));
  INV_X1    g299(.A(G1gat), .ZN(new_n501_));
  INV_X1    g300(.A(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G1gat), .B(G8gat), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n499_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n497_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n497_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(new_n514_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G169gat), .B(G197gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n520_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT10), .B(G99gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534_));
  AND2_X1   g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(KEYINPUT9), .ZN(new_n536_));
  INV_X1    g335(.A(G85gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n536_), .B1(new_n540_), .B2(KEYINPUT9), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n533_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT7), .ZN(new_n543_));
  INV_X1    g342(.A(G99gat), .ZN(new_n544_));
  INV_X1    g343(.A(G106gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(new_n530_), .A3(new_n531_), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT8), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n535_), .A2(new_n534_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n549_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n542_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G71gat), .B(G78gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT11), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n557_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n554_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n562_), .B(new_n542_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT65), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT66), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n554_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n548_), .A2(new_n550_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT8), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n572_), .A2(new_n551_), .B1(new_n533_), .B2(new_n541_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT66), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n570_), .A2(new_n574_), .A3(KEYINPUT12), .A4(new_n563_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n565_), .A2(KEYINPUT12), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n564_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n577_), .A3(new_n567_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n567_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT65), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT67), .ZN(new_n584_));
  XOR2_X1   g383(.A(G176gat), .B(G204gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n568_), .A2(new_n578_), .A3(new_n581_), .A4(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT68), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n579_), .A2(new_n580_), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT65), .B(new_n567_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n592_), .A2(KEYINPUT68), .A3(new_n578_), .A4(new_n586_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n578_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n586_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n594_), .A2(KEYINPUT13), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT13), .B1(new_n594_), .B2(new_n597_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n525_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n597_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(KEYINPUT13), .A3(new_n597_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(KEYINPUT69), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n524_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n490_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n570_), .A2(new_n574_), .A3(new_n499_), .ZN(new_n609_));
  OR2_X1    g408(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n610_));
  NAND2_X1  g409(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(G232gat), .ZN(new_n613_));
  INV_X1    g412(.A(G233gat), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n610_), .B(new_n611_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT35), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT35), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n620_), .A3(new_n617_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT71), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n573_), .B2(new_n511_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n609_), .A2(new_n619_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT72), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n609_), .A2(KEYINPUT72), .A3(new_n623_), .A4(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n609_), .A2(new_n623_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n619_), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n626_), .A2(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G190gat), .B(G218gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(KEYINPUT36), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n608_), .B1(new_n630_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n626_), .A2(new_n627_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n628_), .A2(new_n629_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n633_), .B(KEYINPUT36), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n640_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n639_), .B2(KEYINPUT73), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT73), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n630_), .A2(new_n645_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n644_), .A2(new_n646_), .B1(new_n635_), .B2(new_n630_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n647_), .B2(KEYINPUT37), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n510_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n508_), .A2(G231gat), .A3(G233gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n562_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n563_), .A3(new_n651_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT16), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G183gat), .B(G211gat), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n658_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT17), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n655_), .B1(KEYINPUT76), .B2(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(KEYINPUT76), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n661_), .A2(KEYINPUT17), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT75), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n655_), .A2(KEYINPUT74), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT74), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n653_), .A2(new_n671_), .A3(new_n654_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n666_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n648_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n607_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n501_), .A3(new_n358_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT38), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT99), .Z(new_n680_));
  NOR2_X1   g479(.A1(new_n647_), .A2(new_n674_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n607_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n501_), .B1(new_n683_), .B2(new_n358_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n678_), .B2(new_n677_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n680_), .A2(new_n685_), .ZN(G1324gat));
  NOR2_X1   g485(.A1(new_n486_), .A2(new_n487_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G8gat), .B1(new_n682_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT39), .ZN(new_n689_));
  INV_X1    g488(.A(new_n687_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n676_), .A2(new_n502_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n682_), .B2(new_n478_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n695_), .A2(KEYINPUT41), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(KEYINPUT41), .ZN(new_n697_));
  INV_X1    g496(.A(G15gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n676_), .A2(new_n698_), .A3(new_n477_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n699_), .ZN(G1326gat));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n443_), .B(KEYINPUT101), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n683_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT42), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n676_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1327gat));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n490_), .A2(KEYINPUT103), .A3(new_n707_), .A4(new_n648_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n489_), .A2(new_n485_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n477_), .B1(new_n442_), .B2(new_n451_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n648_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n712_), .B2(KEYINPUT43), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n707_), .B(new_n648_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n708_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n606_), .A2(new_n717_), .A3(new_n674_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n606_), .B2(new_n674_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT104), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n716_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n716_), .B2(new_n720_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(G29gat), .A3(new_n358_), .ZN(new_n726_));
  INV_X1    g525(.A(G29gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n647_), .A2(new_n674_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT105), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n607_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n731_), .B2(new_n444_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n726_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(G1328gat));
  INV_X1    g534(.A(G36gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n730_), .A2(new_n736_), .A3(new_n690_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT45), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n723_), .A2(new_n724_), .A3(new_n687_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n736_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1329gat));
  AOI21_X1  g541(.A(G43gat), .B1(new_n730_), .B2(new_n477_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT108), .ZN(new_n744_));
  INV_X1    g543(.A(G43gat), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n478_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT107), .B1(new_n725_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748_));
  INV_X1    g547(.A(new_n746_), .ZN(new_n749_));
  NOR4_X1   g548(.A1(new_n723_), .A2(new_n724_), .A3(new_n748_), .A4(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n744_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT47), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n753_), .B(new_n744_), .C1(new_n747_), .C2(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1330gat));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n725_), .A2(new_n756_), .A3(new_n443_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G50gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n725_), .B2(new_n443_), .ZN(new_n759_));
  INV_X1    g558(.A(G50gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n702_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT110), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n758_), .A2(new_n759_), .B1(new_n731_), .B2(new_n762_), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n600_), .A2(new_n605_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n490_), .A2(new_n765_), .A3(new_n524_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n681_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n444_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n675_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n769_), .A2(KEYINPUT111), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(KEYINPUT111), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(new_n524_), .A3(new_n490_), .A4(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n358_), .A2(new_n350_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(G1332gat));
  OAI21_X1  g573(.A(G64gat), .B1(new_n767_), .B2(new_n687_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(KEYINPUT48), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(KEYINPUT48), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n687_), .A2(G64gat), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n776_), .A2(new_n777_), .B1(new_n772_), .B2(new_n778_), .ZN(G1333gat));
  OAI21_X1  g578(.A(G71gat), .B1(new_n767_), .B2(new_n478_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT49), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT49), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n478_), .A2(G71gat), .ZN(new_n783_));
  OAI22_X1  g582(.A1(new_n781_), .A2(new_n782_), .B1(new_n772_), .B2(new_n783_), .ZN(G1334gat));
  NAND3_X1  g583(.A1(new_n766_), .A2(new_n681_), .A3(new_n702_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G78gat), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(KEYINPUT50), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(KEYINPUT50), .ZN(new_n788_));
  INV_X1    g587(.A(G78gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n702_), .A2(new_n789_), .ZN(new_n790_));
  OAI22_X1  g589(.A1(new_n787_), .A2(new_n788_), .B1(new_n772_), .B2(new_n790_), .ZN(G1335gat));
  AOI21_X1  g590(.A(new_n668_), .B1(new_n655_), .B2(KEYINPUT74), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n792_), .A2(new_n672_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n523_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n520_), .B(new_n794_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n764_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n716_), .A2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT112), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n537_), .B1(new_n798_), .B2(new_n358_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n766_), .A2(new_n729_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n800_), .A2(G85gat), .A3(new_n444_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1336gat));
  INV_X1    g601(.A(new_n800_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G92gat), .B1(new_n803_), .B2(new_n690_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n687_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT113), .Z(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n798_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n797_), .B2(new_n478_), .ZN(new_n810_));
  OR3_X1    g609(.A1(new_n800_), .A2(new_n526_), .A3(new_n478_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n810_), .A2(new_n811_), .B1(KEYINPUT115), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(KEYINPUT115), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n716_), .A2(new_n796_), .A3(new_n443_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G106gat), .ZN(new_n817_));
  XOR2_X1   g616(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT117), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n816_), .A2(new_n821_), .A3(G106gat), .A4(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n803_), .A2(new_n545_), .A3(new_n443_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT53), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n824_), .A2(new_n828_), .A3(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1339gat));
  NOR2_X1   g629(.A1(new_n690_), .A2(new_n444_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n477_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n630_), .A2(new_n635_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n646_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n640_), .B1(new_n630_), .B2(new_n645_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n837_), .A2(new_n608_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n598_), .A2(new_n599_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT118), .B1(new_n795_), .B2(new_n674_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n524_), .A2(new_n793_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .A4(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n844_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n848_), .A2(KEYINPUT119), .A3(new_n839_), .A4(new_n838_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n840_), .A2(new_n844_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT54), .B1(new_n850_), .B2(new_n648_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n847_), .A2(new_n849_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n644_), .A2(new_n646_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n578_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n575_), .A2(new_n577_), .A3(KEYINPUT55), .A4(new_n567_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n575_), .A2(new_n577_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n567_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(new_n857_), .A3(new_n860_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n861_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT56), .B1(new_n861_), .B2(new_n596_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n795_), .B(new_n594_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n515_), .A2(new_n794_), .A3(new_n518_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n513_), .A2(new_n514_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n867_), .B2(new_n794_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n601_), .A2(new_n868_), .ZN(new_n869_));
  AOI221_X4 g668(.A(new_n853_), .B1(new_n854_), .B2(new_n834_), .C1(new_n864_), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n864_), .A2(new_n869_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n871_), .B2(new_n837_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n594_), .B(new_n868_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n876_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n877_), .A2(new_n648_), .A3(new_n878_), .A4(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n793_), .B1(new_n873_), .B2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n441_), .B(new_n833_), .C1(new_n852_), .C2(new_n881_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n882_), .A2(KEYINPUT59), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n882_), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT121), .B1(new_n882_), .B2(KEYINPUT59), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G113gat), .B1(new_n886_), .B2(new_n524_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n524_), .A2(G113gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n882_), .B2(new_n888_), .ZN(G1340gat));
  OAI21_X1  g688(.A(G120gat), .B1(new_n886_), .B2(new_n764_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n882_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n892_));
  INV_X1    g691(.A(G120gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n765_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n890_), .A2(new_n896_), .ZN(G1341gat));
  INV_X1    g696(.A(G127gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n674_), .A2(new_n898_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n883_), .B(new_n899_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n882_), .B2(new_n674_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT122), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n904_), .A3(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1342gat));
  XOR2_X1   g705(.A(KEYINPUT123), .B(G134gat), .Z(new_n907_));
  NOR3_X1   g706(.A1(new_n886_), .A2(new_n838_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G134gat), .B1(new_n891_), .B2(new_n647_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1343gat));
  NOR2_X1   g709(.A1(new_n852_), .A2(new_n881_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n911_), .A2(new_n477_), .A3(new_n441_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n831_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n524_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n316_), .ZN(G1344gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n764_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n317_), .ZN(G1345gat));
  NOR2_X1   g716(.A1(new_n913_), .A2(new_n674_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT61), .B(G155gat), .Z(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1346gat));
  OAI21_X1  g719(.A(G162gat), .B1(new_n913_), .B2(new_n838_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n837_), .A2(G162gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n913_), .B2(new_n922_), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n687_), .A2(new_n358_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n477_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n911_), .A2(new_n702_), .A3(new_n925_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n926_), .A2(new_n795_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n928_));
  OR3_X1    g727(.A1(new_n927_), .A2(new_n228_), .A3(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n228_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n215_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n930_), .A3(new_n931_), .ZN(G1348gat));
  AOI21_X1  g731(.A(G176gat), .B1(new_n926_), .B2(new_n765_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n911_), .A2(new_n443_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n764_), .A2(new_n216_), .A3(new_n925_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(G1349gat));
  NAND4_X1  g735(.A1(new_n934_), .A2(new_n793_), .A3(new_n477_), .A4(new_n924_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n674_), .A2(new_n236_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n937_), .A2(new_n223_), .B1(new_n926_), .B2(new_n938_), .ZN(G1350gat));
  NAND2_X1  g738(.A1(new_n647_), .A2(new_n240_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT125), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n926_), .A2(new_n941_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n926_), .A2(new_n648_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n224_), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n912_), .A2(new_n924_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n795_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n946_), .A2(new_n949_), .A3(G204gat), .A4(new_n765_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(KEYINPUT126), .B(G204gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n951_), .B1(new_n945_), .B2(new_n764_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n950_), .A2(new_n952_), .ZN(G1353gat));
  NOR2_X1   g752(.A1(new_n945_), .A2(new_n674_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AND2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n957_), .B1(new_n954_), .B2(new_n955_), .ZN(G1354gat));
  AOI21_X1  g757(.A(G218gat), .B1(new_n946_), .B2(new_n647_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n838_), .A2(new_n265_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(KEYINPUT127), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n959_), .B1(new_n946_), .B2(new_n961_), .ZN(G1355gat));
endmodule


