//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT80), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(new_n205_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n206_), .B2(new_n207_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n206_), .A2(new_n207_), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n214_), .A2(new_n216_), .B1(new_n217_), .B2(KEYINPUT3), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n213_), .A2(new_n218_), .A3(KEYINPUT81), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT81), .B1(new_n213_), .B2(new_n218_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n202_), .B(new_n204_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G127gat), .B(G134gat), .Z(new_n222_));
  XOR2_X1   g021(.A(G113gat), .B(G120gat), .Z(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n206_), .A2(new_n207_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n203_), .B1(KEYINPUT1), .B2(new_n202_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n228_));
  AOI211_X1 g027(.A(new_n210_), .B(new_n226_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n221_), .A2(new_n225_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n204_), .A2(new_n202_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n213_), .A2(new_n218_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n213_), .A2(new_n218_), .A3(KEYINPUT81), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n224_), .B1(new_n237_), .B2(new_n229_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n239_));
  OAI211_X1 g038(.A(KEYINPUT4), .B(new_n231_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n221_), .A2(new_n230_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(KEYINPUT86), .A3(new_n244_), .A4(new_n224_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n238_), .A2(new_n231_), .A3(new_n241_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT87), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n238_), .A2(new_n231_), .A3(new_n249_), .A4(new_n241_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G1gat), .B(G29gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G85gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G169gat), .B(G176gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n257_), .B1(new_n259_), .B2(KEYINPUT24), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G183gat), .A3(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT23), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT78), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n263_), .B2(KEYINPUT23), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n262_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT77), .B(G190gat), .Z(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(KEYINPUT26), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT25), .B(G183gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n260_), .B(new_n268_), .C1(new_n271_), .C2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n262_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n261_), .B1(G183gat), .B2(G190gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT79), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n263_), .B2(KEYINPUT23), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n277_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n270_), .A2(G183gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n276_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G43gat), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n274_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n274_), .B2(new_n285_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n224_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(G15gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT30), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT31), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n224_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n290_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n255_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n246_), .A2(new_n299_), .A3(new_n248_), .A4(new_n250_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n256_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G106gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n221_), .B2(new_n230_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G211gat), .B(G218gat), .Z(new_n305_));
  INV_X1    g104(.A(KEYINPUT21), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(KEYINPUT84), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n310_));
  INV_X1    g109(.A(G197gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(G204gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(KEYINPUT21), .A3(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n307_), .A2(new_n306_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n308_), .A2(new_n313_), .B1(new_n305_), .B2(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n304_), .A2(G78gat), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G78gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT29), .B1(new_n237_), .B2(new_n229_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n313_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n305_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n302_), .B1(new_n316_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(G78gat), .B1(new_n304_), .B2(new_n315_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(G106gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G22gat), .B(G50gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n331_));
  OR4_X1    g130(.A1(KEYINPUT28), .A2(new_n237_), .A3(KEYINPUT29), .A4(new_n229_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT28), .B1(new_n243_), .B2(KEYINPUT29), .ZN(new_n333_));
  INV_X1    g132(.A(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n335_), .A2(G228gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(G228gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT83), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n332_), .A2(new_n333_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n342_));
  OAI22_X1  g141(.A1(new_n330_), .A2(new_n331_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT20), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n274_), .A2(new_n285_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(new_n321_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n264_), .A2(KEYINPUT79), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n262_), .B1(new_n349_), .B2(new_n281_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n258_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n272_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n350_), .A2(new_n352_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n278_), .A2(new_n266_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n267_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n277_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n276_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n315_), .A2(new_n357_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n345_), .B1(new_n348_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n354_), .B(new_n356_), .C1(new_n258_), .C2(new_n351_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(new_n283_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n276_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n361_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n268_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n321_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n315_), .A2(new_n274_), .A3(new_n285_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(KEYINPUT20), .A4(new_n345_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT18), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n365_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n373_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n364_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT27), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n345_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT92), .B1(new_n367_), .B2(new_n370_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n362_), .A2(new_n357_), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n315_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n383_), .B1(new_n387_), .B2(new_n348_), .ZN(new_n388_));
  AND4_X1   g187(.A1(KEYINPUT20), .A2(new_n371_), .A3(new_n383_), .A4(new_n372_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n377_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT93), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(KEYINPUT93), .B(new_n377_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n381_), .A2(KEYINPUT27), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n382_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n316_), .A2(new_n322_), .A3(new_n302_), .ZN(new_n397_));
  AOI21_X1  g196(.A(G106gat), .B1(new_n324_), .B2(new_n325_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n327_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n341_), .A2(new_n342_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n329_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n301_), .A2(new_n343_), .A3(new_n396_), .A4(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT95), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n256_), .A2(new_n300_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n399_), .A2(new_n400_), .A3(new_n329_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n400_), .B1(new_n399_), .B2(new_n329_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n405_), .B(new_n396_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n343_), .A2(new_n401_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n411_), .A2(KEYINPUT94), .A3(new_n405_), .A4(new_n396_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n378_), .A2(new_n381_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n240_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT90), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n238_), .A2(new_n231_), .A3(new_n242_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n416_), .A2(new_n255_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n413_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT88), .B1(new_n300_), .B2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n246_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(KEYINPUT33), .A4(new_n299_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT33), .B1(new_n300_), .B2(KEYINPUT89), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(KEYINPUT89), .B2(new_n300_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n256_), .A2(new_n300_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n380_), .A2(new_n364_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n379_), .A2(KEYINPUT32), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n430_), .A2(KEYINPUT91), .A3(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT91), .B1(new_n430_), .B2(new_n432_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n426_), .A2(new_n428_), .B1(new_n429_), .B2(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n410_), .B(new_n412_), .C1(new_n437_), .C2(new_n411_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n298_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n404_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441_));
  INV_X1    g240(.A(G1gat), .ZN(new_n442_));
  INV_X1    g241(.A(G8gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G8gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  XOR2_X1   g246(.A(G29gat), .B(G36gat), .Z(new_n448_));
  XOR2_X1   g247(.A(G43gat), .B(G50gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n448_), .B(new_n449_), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n445_), .B(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT76), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(G229gat), .A3(G233gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n450_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n453_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n451_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G169gat), .B(G197gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n458_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n440_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  AND2_X1   g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT9), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n476_), .A2(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT9), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n481_), .A2(new_n486_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n302_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n477_), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n494_), .B(new_n497_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT65), .B1(new_n479_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n489_), .A2(new_n503_), .A3(new_n490_), .ZN(new_n504_));
  AND4_X1   g303(.A1(new_n493_), .A2(new_n500_), .A3(new_n502_), .A4(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n502_), .A2(new_n504_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n493_), .B1(new_n506_), .B2(new_n500_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n492_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n512_));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513_));
  OR2_X1    g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n513_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n497_), .A2(new_n494_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n502_), .A2(new_n504_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT8), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n506_), .A2(new_n493_), .A3(new_n500_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(KEYINPUT66), .A3(new_n492_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n510_), .A2(new_n518_), .A3(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n505_), .A2(new_n507_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n492_), .A2(KEYINPUT67), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n481_), .A2(new_n486_), .A3(new_n529_), .A4(new_n491_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT68), .B1(new_n527_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT68), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n524_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n518_), .A2(KEYINPUT12), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n474_), .A2(new_n526_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n510_), .A2(new_n525_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n517_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n517_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n526_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n541_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G120gat), .B(G148gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT13), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT13), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT70), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT72), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n536_), .A2(new_n460_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n452_), .B1(new_n510_), .B2(new_n525_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT35), .B(new_n569_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n536_), .A2(new_n460_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n567_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n566_), .B1(new_n578_), .B2(new_n565_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT73), .B1(new_n572_), .B2(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n582_), .B(new_n566_), .C1(new_n578_), .C2(new_n565_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT74), .B(KEYINPUT37), .Z(new_n584_));
  AND3_X1   g383(.A1(new_n581_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n517_), .B(new_n588_), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT75), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n447_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G127gat), .B(G155gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT16), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n590_), .B(new_n453_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n595_), .B(KEYINPUT17), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n587_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n473_), .A2(new_n561_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n442_), .A3(new_n429_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n581_), .A2(new_n583_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT96), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n440_), .A2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n560_), .A2(new_n472_), .A3(new_n602_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n405_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n606_), .A2(new_n607_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n615_), .A3(new_n616_), .ZN(G1324gat));
  INV_X1    g416(.A(new_n396_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n605_), .A2(new_n443_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620_));
  INV_X1    g419(.A(new_n614_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n618_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n620_), .B1(new_n622_), .B2(G8gat), .ZN(new_n623_));
  AOI211_X1 g422(.A(KEYINPUT39), .B(new_n443_), .C1(new_n621_), .C2(new_n618_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n619_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g425(.A1(new_n604_), .A2(G15gat), .A3(new_n439_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G15gat), .B1(new_n614_), .B2(new_n439_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(G1326gat));
  INV_X1    g431(.A(new_n411_), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n604_), .A2(G22gat), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n621_), .A2(new_n411_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT97), .B(KEYINPUT42), .Z(new_n636_));
  AND3_X1   g435(.A1(new_n635_), .A2(G22gat), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n635_), .B2(G22gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n609_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n602_), .ZN(new_n641_));
  NOR4_X1   g440(.A1(new_n440_), .A2(new_n472_), .A3(new_n560_), .A4(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G29gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n429_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  INV_X1    g444(.A(new_n584_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n609_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n581_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n410_), .A2(new_n412_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n425_), .A2(new_n422_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n420_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n428_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n436_), .A2(new_n429_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n411_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n439_), .B1(new_n650_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n404_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n649_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n645_), .B1(new_n658_), .B2(KEYINPUT98), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n660_), .B(KEYINPUT43), .C1(new_n440_), .C2(new_n649_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n560_), .A2(new_n472_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n602_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT44), .B1(new_n662_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n664_), .C1(new_n659_), .C2(new_n661_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n666_), .A2(new_n668_), .A3(new_n405_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n644_), .B1(new_n669_), .B2(new_n643_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(KEYINPUT101), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n662_), .A2(new_n665_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n667_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n665_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n618_), .A4(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G36gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n666_), .A2(new_n668_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n676_), .B1(new_n680_), .B2(new_n618_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT100), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n675_), .A2(new_n618_), .A3(new_n677_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT99), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(G36gat), .A4(new_n678_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n682_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(G36gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n642_), .A2(new_n688_), .A3(new_n618_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT45), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(KEYINPUT45), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n691_), .A2(new_n692_), .B1(KEYINPUT101), .B2(new_n671_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n673_), .B1(new_n687_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n693_), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n672_), .B(new_n695_), .C1(new_n682_), .C2(new_n686_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1329gat));
  XOR2_X1   g496(.A(KEYINPUT102), .B(G43gat), .Z(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n642_), .B2(new_n298_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT103), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n298_), .A2(G43gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n680_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n642_), .A2(new_n704_), .A3(new_n411_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n680_), .A2(KEYINPUT104), .A3(new_n411_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT104), .B1(new_n680_), .B2(new_n411_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1331gat));
  INV_X1    g508(.A(new_n561_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n602_), .A2(new_n471_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n612_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n405_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n440_), .A2(new_n471_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n560_), .A3(new_n603_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n405_), .A2(G57gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n712_), .B2(new_n396_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n396_), .A2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n715_), .B2(new_n720_), .ZN(G1333gat));
  OR3_X1    g520(.A1(new_n715_), .A2(G71gat), .A3(new_n439_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G71gat), .B1(new_n712_), .B2(new_n439_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(KEYINPUT49), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(KEYINPUT49), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(G1334gat));
  OAI21_X1  g525(.A(G78gat), .B1(new_n712_), .B2(new_n633_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT50), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n411_), .A2(new_n317_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n715_), .B2(new_n729_), .ZN(G1335gat));
  NAND4_X1  g529(.A1(new_n714_), .A2(new_n710_), .A3(new_n602_), .A4(new_n640_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n487_), .A3(new_n429_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n560_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n602_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n471_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n662_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n659_), .A2(KEYINPUT105), .A3(new_n661_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n429_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n733_), .B1(new_n742_), .B2(new_n487_), .ZN(G1336gat));
  NAND3_X1  g542(.A1(new_n732_), .A2(new_n488_), .A3(new_n618_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n741_), .A2(new_n618_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n488_), .ZN(G1337gat));
  AOI21_X1  g545(.A(new_n496_), .B1(new_n741_), .B2(new_n298_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n298_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n732_), .B2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g549(.A1(new_n732_), .A2(new_n411_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n737_), .A2(new_n633_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n302_), .B1(new_n662_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n754_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n751_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762_));
  INV_X1    g561(.A(new_n711_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n560_), .B2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n711_), .A2(new_n558_), .A3(KEYINPUT107), .A4(new_n559_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n649_), .A3(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n766_), .B(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n457_), .A2(new_n462_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n462_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n467_), .B1(new_n461_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n470_), .A2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n557_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n471_), .A2(new_n554_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT109), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n471_), .A2(new_n554_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n526_), .A2(new_n474_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n527_), .A2(KEYINPUT68), .A3(new_n531_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n534_), .B1(new_n533_), .B2(new_n524_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n538_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n785_), .A3(new_n545_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n541_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n539_), .B2(new_n543_), .ZN(new_n789_));
  AND4_X1   g588(.A1(new_n788_), .A2(new_n543_), .A3(new_n785_), .A4(new_n782_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT110), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n782_), .A2(new_n785_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n545_), .A2(new_n540_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT55), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n539_), .A2(new_n788_), .A3(new_n543_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n787_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n792_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n552_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n781_), .B1(new_n801_), .B2(KEYINPUT111), .ZN(new_n802_));
  AOI221_X4 g601(.A(KEYINPUT110), .B1(new_n541_), .B2(new_n786_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n798_), .B1(new_n797_), .B2(new_n787_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n552_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n776_), .B1(new_n802_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n770_), .B1(new_n811_), .B2(new_n640_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n776_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n806_), .B(new_n553_), .C1(new_n792_), .C2(new_n799_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n801_), .A2(new_n814_), .A3(KEYINPUT111), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n778_), .A2(new_n780_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n640_), .A2(new_n770_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n812_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n555_), .A2(new_n775_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT58), .B(new_n822_), .C1(new_n801_), .C2(new_n814_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT112), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n807_), .A2(new_n809_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(KEYINPUT58), .A4(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n822_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n649_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n822_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n587_), .B1(new_n836_), .B2(KEYINPUT58), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT113), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n821_), .A2(new_n834_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n769_), .B1(new_n840_), .B2(new_n602_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n633_), .A2(new_n298_), .A3(new_n429_), .A4(new_n396_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n832_), .A2(new_n812_), .A3(new_n820_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n769_), .B1(new_n844_), .B2(new_n602_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT114), .B(KEYINPUT59), .Z(new_n847_));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n842_), .B2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n846_), .B(new_n849_), .C1(new_n848_), .C2(new_n842_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n843_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n472_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n841_), .A2(new_n842_), .ZN(new_n853_));
  INV_X1    g652(.A(G113gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n471_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(G1340gat));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n734_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n853_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n857_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n851_), .A2(new_n561_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT116), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n859_), .C1(new_n860_), .C2(new_n857_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n851_), .B2(new_n602_), .ZN(new_n866_));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n853_), .A2(new_n867_), .A3(new_n735_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1342gat));
  AOI21_X1  g668(.A(G134gat), .B1(new_n853_), .B2(new_n611_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n851_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n587_), .A2(G134gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT117), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n870_), .B1(new_n871_), .B2(new_n873_), .ZN(G1343gat));
  NOR2_X1   g673(.A1(new_n633_), .A2(new_n298_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n618_), .A2(new_n405_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n812_), .A2(new_n820_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT113), .B1(new_n828_), .B2(new_n831_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n735_), .B1(new_n879_), .B2(new_n839_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n875_), .B(new_n876_), .C1(new_n880_), .C2(new_n769_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT118), .ZN(new_n882_));
  INV_X1    g681(.A(new_n875_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n812_), .B(new_n820_), .C1(new_n838_), .C2(KEYINPUT113), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n832_), .A2(new_n833_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n602_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n769_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n883_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n876_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n882_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n471_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT119), .B(G141gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1344gat));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n710_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n891_), .B2(new_n735_), .ZN(new_n900_));
  AOI211_X1 g699(.A(KEYINPUT120), .B(new_n602_), .C1(new_n882_), .C2(new_n890_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n889_), .B1(new_n888_), .B2(new_n876_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n876_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n841_), .A2(KEYINPUT118), .A3(new_n883_), .A4(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n735_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT120), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n891_), .A2(new_n899_), .A3(new_n735_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n897_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n902_), .A2(new_n909_), .ZN(G1346gat));
  AOI21_X1  g709(.A(G162gat), .B1(new_n891_), .B2(new_n611_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n587_), .A2(G162gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT121), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n891_), .B2(new_n913_), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n396_), .A2(new_n429_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n439_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n411_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n471_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n735_), .B1(new_n821_), .B2(new_n832_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT122), .B(new_n921_), .C1(new_n922_), .C2(new_n769_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n845_), .B2(new_n920_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n925_), .A3(G169gat), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n923_), .A2(new_n925_), .A3(KEYINPUT123), .A4(G169gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(KEYINPUT62), .A3(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n926_), .A2(new_n927_), .A3(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT22), .B(G169gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n846_), .A2(new_n921_), .A3(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(new_n932_), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT124), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n930_), .A2(new_n937_), .A3(new_n932_), .A4(new_n934_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1348gat));
  NOR3_X1   g738(.A1(new_n845_), .A2(new_n411_), .A3(new_n918_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n941_), .A2(G176gat), .A3(new_n734_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n841_), .B2(new_n411_), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT125), .B(new_n633_), .C1(new_n880_), .C2(new_n769_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n944_), .A2(new_n945_), .A3(new_n710_), .A4(new_n917_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n942_), .B1(new_n946_), .B2(G176gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(KEYINPUT126), .ZN(G1349gat));
  NAND3_X1  g747(.A1(new_n940_), .A2(new_n273_), .A3(new_n735_), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(KEYINPUT127), .Z(new_n950_));
  NAND4_X1  g749(.A1(new_n944_), .A2(new_n945_), .A3(new_n735_), .A4(new_n917_), .ZN(new_n951_));
  INV_X1    g750(.A(G183gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n941_), .B2(new_n649_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n940_), .A2(new_n353_), .A3(new_n611_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n841_), .A2(new_n883_), .A3(new_n916_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n471_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n710_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g760(.A1(new_n957_), .A2(new_n735_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  AND2_X1   g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n962_), .A2(new_n963_), .A3(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n962_), .B2(new_n963_), .ZN(G1354gat));
  INV_X1    g765(.A(G218gat), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n957_), .A2(new_n967_), .A3(new_n611_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n957_), .A2(new_n587_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n967_), .ZN(G1355gat));
endmodule


