//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n963_, new_n964_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n987_, new_n989_,
    new_n990_, new_n992_, new_n993_, new_n995_, new_n996_, new_n997_,
    new_n999_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_;
  XNOR2_X1  g000(.A(G113gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G120gat), .B(G127gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n203_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(KEYINPUT86), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT86), .ZN(new_n208_));
  INV_X1    g007(.A(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(new_n204_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT87), .B1(new_n215_), .B2(KEYINPUT1), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n214_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n215_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(new_n218_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n211_), .B(KEYINPUT3), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n213_), .B(KEYINPUT2), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n207_), .B(new_n210_), .C1(new_n221_), .C2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n217_), .A2(new_n218_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n216_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n220_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n213_), .A3(new_n212_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n225_), .A2(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n223_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n232_), .B(new_n234_), .C1(new_n209_), .C2(new_n204_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G1gat), .B(G29gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT0), .ZN(new_n239_));
  INV_X1    g038(.A(G57gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G85gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT94), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n228_), .B2(KEYINPUT4), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n207_), .A2(new_n210_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n232_), .A2(new_n234_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n245_), .A2(KEYINPUT94), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n228_), .A2(new_n235_), .A3(KEYINPUT4), .ZN(new_n250_));
  INV_X1    g049(.A(new_n236_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n237_), .B(new_n242_), .C1(new_n249_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT95), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT33), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT33), .B1(new_n253_), .B2(new_n254_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G169gat), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT82), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT23), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(KEYINPUT82), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n269_), .A2(KEYINPUT92), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(KEYINPUT92), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n258_), .B(new_n261_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G197gat), .B(G204gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(KEYINPUT21), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G190gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT25), .B(G183gat), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G169gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n260_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT24), .A3(new_n258_), .ZN(new_n283_));
  OR3_X1    g082(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(new_n267_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n280_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n272_), .A2(new_n277_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT93), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n272_), .A2(KEYINPUT93), .A3(new_n277_), .A4(new_n289_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n259_), .A2(KEYINPUT84), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n281_), .A2(KEYINPUT22), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n260_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI221_X1 g096(.A(new_n258_), .B1(new_n294_), .B2(new_n297_), .C1(new_n265_), .C2(new_n287_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n264_), .A2(new_n268_), .A3(new_n284_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n283_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n264_), .A2(KEYINPUT83), .A3(new_n268_), .A4(new_n284_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306_));
  INV_X1    g105(.A(G183gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT25), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(KEYINPUT25), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n278_), .B(new_n308_), .C1(new_n309_), .C2(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n283_), .A2(new_n303_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n304_), .A2(new_n305_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n298_), .B1(new_n302_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n277_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n292_), .A2(KEYINPUT20), .A3(new_n293_), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT19), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n261_), .A2(new_n258_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n269_), .A2(KEYINPUT92), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n269_), .A2(KEYINPUT92), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n314_), .B1(new_n324_), .B2(new_n288_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n310_), .A2(new_n311_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n326_), .A2(new_n301_), .A3(new_n305_), .A4(new_n304_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(new_n277_), .A3(new_n298_), .ZN(new_n328_));
  AND4_X1   g127(.A1(KEYINPUT20), .A2(new_n325_), .A3(new_n318_), .A4(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G64gat), .ZN(new_n334_));
  INV_X1    g133(.A(G92gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n329_), .B1(new_n319_), .B2(new_n316_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n336_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n244_), .A2(new_n248_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n236_), .A3(new_n250_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n242_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n228_), .A2(new_n235_), .A3(new_n251_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n337_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT96), .B1(new_n257_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n253_), .A2(new_n254_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT33), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT33), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n320_), .A2(new_n330_), .A3(new_n339_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n339_), .B1(new_n320_), .B2(new_n330_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n352_), .A2(new_n355_), .A3(new_n356_), .A4(new_n345_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n325_), .A2(KEYINPUT20), .A3(new_n319_), .A4(new_n328_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n358_), .A2(KEYINPUT99), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(KEYINPUT99), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n315_), .A2(new_n290_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n318_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT98), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(KEYINPUT98), .A3(new_n318_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(KEYINPUT32), .A3(new_n336_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n237_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n250_), .A2(new_n251_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n341_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT100), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n242_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n374_), .B1(new_n373_), .B2(new_n242_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n253_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n331_), .B1(new_n378_), .B2(new_n339_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n370_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n347_), .A2(new_n357_), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n232_), .A2(new_n234_), .A3(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n221_), .A2(new_n227_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n385_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n386_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT91), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n387_), .B2(new_n383_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n247_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(G228gat), .A2(G233gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n277_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n403_));
  OAI21_X1  g202(.A(new_n314_), .B1(new_n387_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n400_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n382_), .B1(new_n395_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n393_), .A2(new_n394_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n394_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n391_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n409_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n382_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n399_), .A2(new_n401_), .B1(new_n404_), .B2(new_n400_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n407_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n410_), .B1(new_n407_), .B2(new_n416_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n313_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n327_), .A2(KEYINPUT30), .A3(new_n298_), .ZN(new_n422_));
  INV_X1    g221(.A(G227gat), .ZN(new_n423_));
  INV_X1    g222(.A(G233gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n421_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G71gat), .B(G99gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n421_), .A2(new_n422_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n425_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n430_), .B1(new_n434_), .B2(new_n427_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G43gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT31), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n207_), .A2(new_n210_), .A3(new_n438_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT85), .B1(new_n444_), .B2(new_n439_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n437_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n437_), .ZN(new_n447_));
  OAI22_X1  g246(.A1(new_n432_), .A2(new_n435_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n446_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n434_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n431_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n419_), .A2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n452_), .B(new_n448_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n395_), .A2(new_n406_), .A3(new_n382_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n414_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n458_));
  OAI22_X1  g257(.A1(new_n457_), .A2(new_n458_), .B1(new_n409_), .B2(new_n408_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n407_), .A2(new_n416_), .A3(new_n410_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n377_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT27), .B1(new_n337_), .B2(new_n340_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n336_), .B1(new_n361_), .B2(new_n368_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT101), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT27), .B1(new_n338_), .B2(new_n339_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n463_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n381_), .A2(new_n455_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n474_), .A2(new_n477_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT8), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n480_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G71gat), .B(G78gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT11), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n240_), .A2(G64gat), .ZN(new_n492_));
  INV_X1    g291(.A(G64gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(G57gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n491_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(G57gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n240_), .A2(G64gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT11), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n490_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n490_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT64), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT10), .B(G99gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(G106gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(KEYINPUT64), .A3(new_n473_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n481_), .A2(new_n482_), .A3(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(G85gat), .A3(G92gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n477_), .A2(new_n513_), .A3(new_n478_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n489_), .A2(new_n502_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT69), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT66), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT64), .B1(new_n508_), .B2(new_n473_), .ZN(new_n525_));
  NOR4_X1   g324(.A1(new_n506_), .A2(new_n507_), .A3(new_n503_), .A4(G106gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n512_), .A2(new_n514_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n510_), .A2(new_n515_), .A3(KEYINPUT66), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n489_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT67), .B1(new_n499_), .B2(new_n501_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n490_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT11), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT11), .B1(new_n496_), .B2(new_n497_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n500_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n532_), .B1(new_n533_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n489_), .A2(new_n516_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n502_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n541_), .A2(KEYINPUT68), .B1(new_n544_), .B2(new_n532_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n531_), .A2(new_n540_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n523_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n517_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n518_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G120gat), .B(G148gat), .ZN(new_n552_));
  INV_X1    g351(.A(G204gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT5), .B(G176gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT70), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n548_), .A2(new_n551_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT13), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G169gat), .ZN(new_n568_));
  INV_X1    g367(.A(G197gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT78), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT75), .B(G1gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(G8gat), .ZN(new_n573_));
  INV_X1    g372(.A(G8gat), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT75), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(G1gat), .ZN(new_n576_));
  INV_X1    g375(.A(G1gat), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(KEYINPUT75), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n574_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT72), .B(G1gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT73), .B(G8gat), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT14), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n577_), .A2(KEYINPUT72), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(G1gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n574_), .A2(KEYINPUT73), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(G8gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n586_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G15gat), .B(G22gat), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n581_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  AOI211_X1 g399(.A(new_n598_), .B(new_n580_), .C1(new_n586_), .C2(new_n596_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G29gat), .B(G36gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G43gat), .B(G50gat), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G43gat), .B(G50gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n600_), .A2(new_n601_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT74), .B1(new_n595_), .B2(KEYINPUT14), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT14), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n585_), .B(new_n612_), .C1(new_n590_), .C2(new_n594_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n599_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n580_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n597_), .A2(new_n599_), .A3(new_n581_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n608_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n571_), .B1(new_n610_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n609_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n615_), .A2(new_n616_), .A3(new_n608_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(KEYINPUT78), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n615_), .A2(new_n616_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT15), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n608_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n605_), .A2(KEYINPUT15), .A3(new_n607_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT79), .B1(new_n625_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n632_), .B(new_n629_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n619_), .B(new_n622_), .C1(new_n631_), .C2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n570_), .B1(new_n624_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n624_), .A2(new_n634_), .A3(new_n570_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n566_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n470_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n542_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT35), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT71), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT34), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n641_), .A2(new_n608_), .B1(new_n642_), .B2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n642_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n531_), .A2(new_n630_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n648_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G134gat), .B(G162gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NOR4_X1   g454(.A1(new_n651_), .A2(new_n652_), .A3(KEYINPUT36), .A4(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n655_), .B(KEYINPUT36), .Z(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n652_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n650_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n656_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT37), .ZN(new_n662_));
  NAND2_X1  g461(.A1(G231gat), .A2(G233gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n625_), .B(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n543_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n664_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n502_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(G183gat), .B(G211gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G127gat), .B(G155gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT17), .Z(new_n673_));
  NAND3_X1  g472(.A1(new_n665_), .A2(new_n667_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n533_), .A2(new_n539_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n666_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n664_), .A2(new_n533_), .A3(new_n539_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n672_), .A2(KEYINPUT17), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT77), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n674_), .A2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n662_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n640_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n582_), .A3(new_n377_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n381_), .A2(new_n455_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n462_), .A2(new_n469_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n661_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n681_), .A3(new_n639_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n577_), .B1(new_n693_), .B2(new_n377_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n687_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n686_), .B2(new_n685_), .ZN(G1324gat));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n639_), .A2(new_n681_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n469_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n690_), .A2(new_n699_), .A3(new_n691_), .A4(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n574_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n470_), .A2(new_n661_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(KEYINPUT102), .A3(new_n700_), .A4(new_n699_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT39), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT39), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n708_), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n700_), .A2(new_n583_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n683_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n698_), .B1(new_n710_), .B2(new_n713_), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT103), .B(new_n712_), .C1(new_n707_), .C2(new_n709_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n697_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n709_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n708_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT103), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n710_), .A2(new_n698_), .A3(new_n713_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(KEYINPUT40), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n722_), .ZN(G1325gat));
  INV_X1    g522(.A(G15gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n693_), .B2(new_n454_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT41), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n684_), .A2(new_n724_), .A3(new_n454_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1326gat));
  INV_X1    g527(.A(G22gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n693_), .B2(new_n419_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n684_), .A2(new_n729_), .A3(new_n419_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT104), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(new_n736_), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1327gat));
  NAND2_X1  g537(.A1(new_n681_), .A2(new_n661_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT106), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n640_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G29gat), .B1(new_n742_), .B2(new_n377_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n662_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n745_), .B2(KEYINPUT105), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n747_), .B(new_n748_), .C1(new_n470_), .C2(new_n744_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n681_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n639_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n746_), .A2(new_n749_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n746_), .A2(KEYINPUT44), .A3(new_n749_), .A4(new_n751_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n377_), .A2(G29gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n743_), .B1(new_n756_), .B2(new_n757_), .ZN(G1328gat));
  NOR2_X1   g557(.A1(new_n469_), .A2(G36gat), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n742_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n760_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n759_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n741_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n754_), .A2(new_n700_), .A3(new_n755_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G36gat), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n768_), .A2(new_n769_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n767_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n770_), .A2(new_n773_), .ZN(G1329gat));
  INV_X1    g573(.A(G43gat), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n453_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n754_), .A2(new_n755_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n754_), .A2(KEYINPUT109), .A3(new_n755_), .A4(new_n776_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n775_), .B1(new_n741_), .B2(new_n453_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT47), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n779_), .A2(new_n784_), .A3(new_n780_), .A4(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1330gat));
  AOI21_X1  g585(.A(G50gat), .B1(new_n742_), .B2(new_n419_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n419_), .A2(G50gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n756_), .B2(new_n788_), .ZN(G1331gat));
  INV_X1    g588(.A(new_n377_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT110), .B1(new_n470_), .B2(new_n638_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n792_));
  INV_X1    g591(.A(new_n638_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n690_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n791_), .A2(new_n794_), .A3(new_n682_), .A4(new_n565_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n790_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n796_), .B2(new_n795_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n793_), .A2(new_n750_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n692_), .A2(new_n566_), .A3(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n790_), .A2(new_n240_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n798_), .A2(new_n240_), .B1(new_n800_), .B2(new_n801_), .ZN(G1332gat));
  AOI21_X1  g601(.A(new_n493_), .B1(new_n800_), .B2(new_n700_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT48), .Z(new_n804_));
  NAND2_X1  g603(.A1(new_n700_), .A2(new_n493_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT112), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n795_), .B2(new_n806_), .ZN(G1333gat));
  INV_X1    g606(.A(G71gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n800_), .B2(new_n454_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT49), .Z(new_n810_));
  NAND2_X1  g609(.A1(new_n454_), .A2(new_n808_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n795_), .B2(new_n811_), .ZN(G1334gat));
  INV_X1    g611(.A(G78gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n800_), .B2(new_n419_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n419_), .A2(new_n813_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n795_), .B2(new_n817_), .ZN(G1335gat));
  NAND4_X1  g617(.A1(new_n791_), .A2(new_n794_), .A3(new_n565_), .A4(new_n740_), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n819_), .A2(G85gat), .A3(new_n790_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n566_), .A2(new_n750_), .A3(new_n638_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n746_), .A2(new_n749_), .A3(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G85gat), .B1(new_n822_), .B2(new_n790_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1336gat));
  OAI21_X1  g623(.A(G92gat), .B1(new_n822_), .B2(new_n469_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n700_), .A2(new_n335_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n819_), .B2(new_n826_), .ZN(G1337gat));
  OAI21_X1  g626(.A(G99gat), .B1(new_n822_), .B2(new_n453_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n454_), .A2(new_n508_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n828_), .B(KEYINPUT114), .C1(new_n819_), .C2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n746_), .A2(new_n419_), .A3(new_n749_), .A4(new_n821_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G106gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n833_), .A2(new_n834_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n832_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n473_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(KEYINPUT52), .C1(new_n834_), .C2(new_n833_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n419_), .A2(new_n473_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n819_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(new_n840_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT53), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n838_), .A2(new_n844_), .A3(new_n840_), .A4(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1339gat));
  INV_X1    g648(.A(G113gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n469_), .A2(new_n377_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n456_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n618_), .A2(new_n619_), .A3(new_n623_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n570_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n622_), .A2(new_n620_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n548_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n637_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n637_), .A2(new_n858_), .A3(KEYINPUT119), .A4(new_n859_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n541_), .A2(KEYINPUT68), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n544_), .A2(new_n532_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n547_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n522_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n521_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n865_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n523_), .A2(new_n545_), .A3(KEYINPUT55), .A4(new_n547_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n866_), .A2(new_n517_), .A3(new_n547_), .A4(new_n867_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n550_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(new_n873_), .A3(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(KEYINPUT56), .A3(new_n557_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n876_), .B2(new_n557_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n853_), .B1(new_n864_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n862_), .A2(new_n863_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(KEYINPUT58), .C1(new_n879_), .C2(new_n878_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n881_), .A2(KEYINPUT120), .A3(new_n662_), .A4(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n637_), .A2(new_n858_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n561_), .A2(new_n886_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n624_), .A2(new_n634_), .A3(new_n570_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n859_), .B1(new_n888_), .B2(new_n635_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(KEYINPUT118), .B2(new_n879_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n876_), .A2(new_n557_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n877_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n887_), .B1(new_n890_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n885_), .B1(new_n896_), .B2(new_n661_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n884_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n881_), .A2(new_n662_), .A3(new_n883_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n890_), .A2(new_n895_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n887_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n661_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n899_), .A2(new_n900_), .B1(new_n903_), .B2(KEYINPUT57), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n750_), .B1(new_n898_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n566_), .A2(new_n907_), .A3(new_n750_), .A4(new_n793_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT117), .B1(new_n799_), .B2(new_n565_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n906_), .B1(new_n910_), .B2(new_n744_), .ZN(new_n911_));
  AOI211_X1 g710(.A(KEYINPUT54), .B(new_n662_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n852_), .B1(new_n905_), .B2(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n850_), .B1(new_n914_), .B2(new_n793_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT121), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n852_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n744_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(KEYINPUT54), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n910_), .A2(new_n906_), .A3(new_n744_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n901_), .A2(new_n902_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(KEYINPUT57), .A3(new_n691_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(new_n897_), .A3(new_n899_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n681_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n918_), .B1(new_n922_), .B2(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n914_), .B2(KEYINPUT59), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n929_), .A2(new_n850_), .A3(new_n793_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n916_), .A2(new_n930_), .ZN(G1340gat));
  INV_X1    g730(.A(new_n852_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n899_), .A2(new_n900_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n933_), .A2(new_n897_), .A3(new_n884_), .A4(new_n924_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n681_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n932_), .B1(new_n935_), .B2(new_n922_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n566_), .A2(G120gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(KEYINPUT60), .B2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n938_), .A2(new_n928_), .A3(new_n565_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(G120gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n940_), .B1(KEYINPUT60), .B2(new_n938_), .ZN(G1341gat));
  OAI21_X1  g740(.A(G127gat), .B1(new_n929_), .B2(new_n681_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n681_), .A2(G127gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n914_), .B2(new_n943_), .ZN(G1342gat));
  INV_X1    g743(.A(G134gat), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n945_), .B1(new_n928_), .B2(new_n662_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n914_), .A2(G134gat), .A3(new_n691_), .ZN(new_n947_));
  OAI21_X1  g746(.A(KEYINPUT122), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n925_), .A2(new_n681_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n917_), .B(new_n852_), .C1(new_n949_), .C2(new_n913_), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n662_), .B(new_n950_), .C1(new_n936_), .C2(new_n917_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(G134gat), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953_));
  INV_X1    g752(.A(new_n947_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n952_), .A2(new_n953_), .A3(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n948_), .A2(new_n955_), .ZN(G1343gat));
  NOR2_X1   g755(.A1(new_n905_), .A2(new_n913_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n957_), .A2(new_n461_), .A3(new_n851_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n638_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n565_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g761(.A1(new_n958_), .A2(new_n750_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT61), .B(G155gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1346gat));
  INV_X1    g764(.A(new_n958_), .ZN(new_n966_));
  OAI21_X1  g765(.A(G162gat), .B1(new_n966_), .B2(new_n744_), .ZN(new_n967_));
  INV_X1    g766(.A(G162gat), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n958_), .A2(new_n968_), .A3(new_n661_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n967_), .A2(new_n969_), .ZN(G1347gat));
  XNOR2_X1  g769(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n971_));
  INV_X1    g770(.A(new_n971_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n949_), .A2(new_n913_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n469_), .A2(new_n377_), .ZN(new_n974_));
  INV_X1    g773(.A(new_n974_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n975_), .A2(new_n453_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n976_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n977_));
  OR2_X1    g776(.A1(new_n973_), .A2(new_n977_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n978_), .A2(new_n793_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n972_), .B1(new_n979_), .B2(new_n281_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n259_), .ZN(new_n981_));
  OAI211_X1 g780(.A(G169gat), .B(new_n971_), .C1(new_n978_), .C2(new_n793_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n980_), .A2(new_n981_), .A3(new_n982_), .ZN(G1348gat));
  INV_X1    g782(.A(new_n978_), .ZN(new_n984_));
  AOI21_X1  g783(.A(G176gat), .B1(new_n984_), .B2(new_n565_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n957_), .A2(new_n419_), .ZN(new_n986_));
  NOR4_X1   g785(.A1(new_n975_), .A2(new_n260_), .A3(new_n453_), .A4(new_n566_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n985_), .B1(new_n986_), .B2(new_n987_), .ZN(G1349gat));
  NOR3_X1   g787(.A1(new_n978_), .A2(new_n681_), .A3(new_n279_), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n986_), .A2(new_n750_), .A3(new_n976_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n989_), .B1(new_n307_), .B2(new_n990_), .ZN(G1350gat));
  OAI21_X1  g790(.A(G190gat), .B1(new_n978_), .B2(new_n744_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n661_), .A2(new_n278_), .ZN(new_n993_));
  OAI21_X1  g792(.A(new_n992_), .B1(new_n978_), .B2(new_n993_), .ZN(G1351gat));
  INV_X1    g793(.A(new_n461_), .ZN(new_n995_));
  OAI211_X1 g794(.A(new_n995_), .B(new_n974_), .C1(new_n905_), .C2(new_n913_), .ZN(new_n996_));
  NOR2_X1   g795(.A1(new_n996_), .A2(new_n793_), .ZN(new_n997_));
  XNOR2_X1  g796(.A(new_n997_), .B(new_n569_), .ZN(G1352gat));
  NOR2_X1   g797(.A1(new_n996_), .A2(new_n566_), .ZN(new_n999_));
  XNOR2_X1  g798(.A(new_n999_), .B(new_n553_), .ZN(G1353gat));
  NOR2_X1   g799(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1001_));
  AND2_X1   g800(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1002_));
  NOR4_X1   g801(.A1(new_n996_), .A2(new_n681_), .A3(new_n1001_), .A4(new_n1002_), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n1001_), .B1(new_n996_), .B2(new_n681_), .ZN(new_n1004_));
  OR2_X1    g803(.A1(new_n1004_), .A2(KEYINPUT124), .ZN(new_n1005_));
  NAND2_X1  g804(.A1(new_n1004_), .A2(KEYINPUT124), .ZN(new_n1006_));
  AOI21_X1  g805(.A(new_n1003_), .B1(new_n1005_), .B2(new_n1006_), .ZN(G1354gat));
  NOR2_X1   g806(.A1(new_n996_), .A2(new_n691_), .ZN(new_n1008_));
  XNOR2_X1  g807(.A(KEYINPUT125), .B(G218gat), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n662_), .A2(new_n1009_), .ZN(new_n1010_));
  XNOR2_X1  g809(.A(new_n1010_), .B(KEYINPUT126), .ZN(new_n1011_));
  OAI22_X1  g810(.A1(new_n1008_), .A2(new_n1009_), .B1(new_n996_), .B2(new_n1011_), .ZN(new_n1012_));
  NAND2_X1  g811(.A1(new_n1012_), .A2(KEYINPUT127), .ZN(new_n1013_));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014_));
  OAI221_X1 g813(.A(new_n1014_), .B1(new_n996_), .B2(new_n1011_), .C1(new_n1008_), .C2(new_n1009_), .ZN(new_n1015_));
  NAND2_X1  g814(.A1(new_n1013_), .A2(new_n1015_), .ZN(G1355gat));
endmodule


