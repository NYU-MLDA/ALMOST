//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT68), .ZN(new_n203_));
  XOR2_X1   g002(.A(G134gat), .B(G162gat), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n207_));
  XOR2_X1   g006(.A(G29gat), .B(G36gat), .Z(new_n208_));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G29gat), .B(G36gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n217_), .B(new_n220_), .C1(new_n222_), .C2(KEYINPUT64), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n220_), .A2(new_n224_), .A3(KEYINPUT9), .A4(new_n221_), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n216_), .A2(new_n223_), .A3(new_n225_), .A4(new_n229_), .ZN(new_n230_));
  OR3_X1    g029(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT6), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n231_), .B(new_n232_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n220_), .A2(new_n221_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n214_), .B(new_n230_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G232gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT34), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT35), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n230_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n238_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT8), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n247_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT15), .B1(new_n210_), .B2(new_n213_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n210_), .A2(KEYINPUT15), .A3(new_n213_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n241_), .B(new_n246_), .C1(new_n251_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT67), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n230_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n210_), .A2(KEYINPUT15), .A3(new_n213_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(new_n252_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n241_), .A4(new_n246_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n244_), .A2(new_n245_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n257_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT36), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n207_), .B1(new_n268_), .B2(new_n206_), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT69), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n257_), .A2(new_n263_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n264_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n257_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT36), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n205_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n270_), .A3(new_n207_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(KEYINPUT71), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n281_), .A3(new_n279_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(KEYINPUT70), .A2(new_n280_), .B1(new_n282_), .B2(KEYINPUT37), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n280_), .A2(KEYINPUT70), .A3(KEYINPUT37), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n288_));
  XOR2_X1   g087(.A(G71gat), .B(G78gat), .Z(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G15gat), .B(G22gat), .ZN(new_n292_));
  INV_X1    g091(.A(G1gat), .ZN(new_n293_));
  INV_X1    g092(.A(G8gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  XOR2_X1   g097(.A(new_n291_), .B(new_n298_), .Z(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT17), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G155gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT16), .ZN(new_n304_));
  XOR2_X1   g103(.A(G183gat), .B(G211gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n301_), .A2(new_n302_), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(KEYINPUT17), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n301_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n285_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n258_), .B(new_n291_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(KEYINPUT12), .ZN(new_n315_));
  OR3_X1    g114(.A1(new_n251_), .A2(KEYINPUT12), .A3(new_n291_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n314_), .B1(new_n317_), .B2(new_n313_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G120gat), .B(G148gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT5), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n324_), .B(KEYINPUT66), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n318_), .A2(new_n323_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT65), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT13), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n326_), .A2(KEYINPUT13), .A3(new_n328_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n311_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G127gat), .B(G134gat), .Z(new_n337_));
  XOR2_X1   g136(.A(G113gat), .B(G120gat), .Z(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT75), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n339_), .B1(new_n344_), .B2(KEYINPUT75), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT31), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT74), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(G15gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT30), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n347_), .B(new_n350_), .Z(new_n351_));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT24), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n355_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT25), .B(G183gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT26), .B(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n366_), .A3(new_n359_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G169gat), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n362_), .A2(new_n365_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(G43gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n370_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n351_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  OR2_X1    g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G141gat), .A2(G148gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383_));
  INV_X1    g182(.A(G141gat), .ZN(new_n384_));
  INV_X1    g183(.A(G148gat), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .A4(KEYINPUT77), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n387_));
  OAI22_X1  g186(.A1(new_n387_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n379_), .B1(new_n382_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n378_), .A2(KEYINPUT1), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G155gat), .A3(G162gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n393_), .A3(new_n377_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G141gat), .B(G148gat), .Z(new_n395_));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n390_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n345_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n344_), .B(new_n390_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n376_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT4), .B1(new_n345_), .B2(new_n399_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(KEYINPUT94), .Z(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G85gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT0), .B(G57gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n400_), .A2(new_n401_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n406_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n402_), .A2(new_n414_), .A3(new_n403_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n419_), .A3(KEYINPUT98), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT98), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n411_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n375_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n399_), .A2(KEYINPUT29), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT21), .ZN(new_n429_));
  AND2_X1   g228(.A1(G197gat), .A2(G204gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT79), .B(new_n429_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(G197gat), .A2(G204gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G197gat), .A2(G204gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(KEYINPUT21), .A3(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G211gat), .B(G218gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n434_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT79), .B1(new_n438_), .B2(new_n429_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT80), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G218gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G211gat), .ZN(new_n442_));
  INV_X1    g241(.A(G211gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G218gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n430_), .A2(new_n431_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(KEYINPUT21), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT79), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n446_), .B2(KEYINPUT21), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n447_), .A2(new_n449_), .A3(new_n450_), .A4(new_n432_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n445_), .A2(new_n446_), .A3(KEYINPUT81), .A4(KEYINPUT21), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n440_), .A2(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G228gat), .ZN(new_n456_));
  INV_X1    g255(.A(G233gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n428_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n453_), .A2(new_n454_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n450_), .B1(new_n462_), .B2(new_n449_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT80), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT82), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n455_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n428_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n458_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n460_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI221_X4 g270(.A(KEYINPUT82), .B1(new_n454_), .B2(new_n453_), .C1(new_n440_), .C2(new_n451_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n440_), .A2(new_n451_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n473_), .B2(new_n461_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n427_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(KEYINPUT83), .A3(new_n458_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n459_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n426_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(KEYINPUT84), .B(new_n459_), .C1(new_n471_), .C2(new_n476_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT85), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n399_), .A2(KEYINPUT29), .ZN(new_n482_));
  XOR2_X1   g281(.A(G22gat), .B(G50gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT78), .B(KEYINPUT28), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n426_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n459_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n475_), .A2(KEYINPUT83), .A3(new_n458_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT83), .B1(new_n475_), .B2(new_n458_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n487_), .B(new_n488_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT86), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n471_), .A2(new_n476_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n487_), .A4(new_n488_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n486_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT84), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n477_), .A2(new_n478_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .A4(new_n426_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n481_), .A2(new_n496_), .A3(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n477_), .A2(new_n487_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n491_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n486_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT93), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G8gat), .B(G36gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G64gat), .B(G92gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT19), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n367_), .A2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n358_), .A2(new_n366_), .A3(KEYINPUT90), .A4(new_n359_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G176gat), .ZN(new_n518_));
  INV_X1    g317(.A(G169gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT22), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT22), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(G169gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n518_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n517_), .A2(new_n526_), .A3(new_n352_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n352_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n520_), .A2(new_n522_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT89), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n530_), .B1(new_n534_), .B2(new_n518_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(KEYINPUT91), .A3(new_n517_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n364_), .B(KEYINPUT88), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n363_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n529_), .A2(new_n536_), .B1(new_n362_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n513_), .B1(new_n540_), .B2(new_n455_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n542_));
  INV_X1    g341(.A(new_n370_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n465_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n473_), .A2(new_n461_), .A3(new_n370_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT20), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT87), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n363_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n362_), .B1(new_n537_), .B2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT91), .B1(new_n535_), .B2(new_n517_), .ZN(new_n551_));
  AND4_X1   g350(.A1(KEYINPUT91), .A2(new_n517_), .A3(new_n352_), .A4(new_n526_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n465_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  AOI221_X4 g355(.A(new_n511_), .B1(new_n541_), .B2(new_n544_), .C1(new_n556_), .C2(new_n513_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n509_), .B(new_n510_), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n513_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n541_), .A2(new_n544_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT27), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n550_), .A2(new_n527_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n550_), .A2(KEYINPUT96), .A3(new_n527_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n466_), .A2(new_n468_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n544_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n513_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n513_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n548_), .A2(new_n554_), .A3(new_n572_), .A4(new_n555_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n564_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n564_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n511_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n557_), .A2(new_n563_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n562_), .A2(new_n563_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n425_), .A2(new_n502_), .A3(new_n505_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n558_), .A2(KEYINPUT32), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n559_), .A2(new_n580_), .A3(new_n560_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n420_), .A2(new_n581_), .A3(new_n422_), .ZN(new_n582_));
  OAI211_X1 g381(.A(KEYINPUT32), .B(new_n558_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n557_), .A2(new_n561_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT33), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n419_), .A2(new_n586_), .ZN(new_n587_));
  OAI221_X1 g386(.A(new_n411_), .B1(new_n585_), .B2(KEYINPUT33), .C1(new_n417_), .C2(new_n418_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n414_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n589_), .B(new_n412_), .C1(new_n414_), .C2(new_n413_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n587_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n582_), .A2(new_n583_), .B1(new_n584_), .B2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n502_), .A2(new_n505_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n375_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n505_), .A2(new_n502_), .B1(new_n578_), .B2(new_n423_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n579_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n298_), .A2(new_n214_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT72), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n298_), .B2(new_n255_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n298_), .A2(new_n214_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT73), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n608_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT73), .B(new_n611_), .C1(new_n602_), .C2(new_n604_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n596_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n336_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT99), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n293_), .A3(new_n424_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n334_), .A2(new_n613_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n310_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n278_), .A2(new_n270_), .A3(new_n207_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n270_), .B1(new_n278_), .B2(new_n207_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT100), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(KEYINPUT100), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n596_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n621_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n423_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n617_), .A2(new_n618_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n619_), .A2(new_n631_), .A3(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(new_n578_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n294_), .B1(new_n629_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT39), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n616_), .A2(new_n294_), .A3(new_n634_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(G1325gat));
  INV_X1    g439(.A(new_n375_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n629_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G15gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  OR3_X1    g444(.A1(new_n615_), .A2(G15gat), .A3(new_n375_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1326gat));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n502_), .A2(new_n505_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n629_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT42), .Z(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n650_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n615_), .B2(new_n654_), .ZN(G1327gat));
  AND4_X1   g454(.A1(new_n614_), .A2(new_n334_), .A3(new_n310_), .A4(new_n624_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n424_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n596_), .A2(new_n659_), .A3(new_n285_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n280_), .A2(KEYINPUT70), .A3(KEYINPUT37), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n281_), .B1(new_n624_), .B2(KEYINPUT71), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT37), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n624_), .B2(new_n281_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT102), .B(new_n664_), .C1(new_n665_), .C2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n596_), .A2(new_n663_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT43), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n661_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n620_), .A2(new_n309_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n658_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n669_), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT103), .B1(new_n669_), .B2(KEYINPUT43), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n660_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n675_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n424_), .A2(G29gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n657_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n656_), .A2(new_n686_), .A3(new_n634_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT45), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n677_), .A2(new_n634_), .A3(new_n681_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT104), .B1(new_n689_), .B2(G36gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT46), .B(new_n688_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1329gat));
  NAND2_X1  g495(.A1(new_n656_), .A2(new_n641_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(G43gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT106), .Z(new_n700_));
  AND4_X1   g499(.A1(G43gat), .A2(new_n677_), .A3(new_n641_), .A4(new_n681_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(G1330gat));
  INV_X1    g503(.A(G50gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n656_), .A2(new_n705_), .A3(new_n651_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n677_), .A2(new_n651_), .A3(new_n681_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT107), .B1(new_n707_), .B2(G50gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT108), .B(new_n706_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1331gat));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715_));
  INV_X1    g514(.A(new_n311_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(new_n334_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n613_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n596_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n311_), .A2(KEYINPUT109), .A3(new_n333_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT110), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n423_), .B1(new_n721_), .B2(KEYINPUT110), .ZN(new_n723_));
  AOI21_X1  g522(.A(G57gat), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND4_X1   g523(.A1(new_n718_), .A2(new_n628_), .A3(new_n333_), .A4(new_n309_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n424_), .A2(G57gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT111), .ZN(G1332gat));
  INV_X1    g527(.A(G64gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n725_), .B2(new_n634_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT48), .Z(new_n731_));
  INV_X1    g530(.A(new_n721_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n729_), .A3(new_n634_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n725_), .B2(new_n641_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n641_), .A2(new_n735_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT113), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n721_), .B2(new_n740_), .ZN(G1334gat));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n725_), .B2(new_n651_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT50), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n732_), .A2(new_n742_), .A3(new_n651_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  AND4_X1   g545(.A1(new_n333_), .A2(new_n719_), .A3(new_n310_), .A4(new_n624_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n218_), .A3(new_n424_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n333_), .A2(new_n718_), .A3(new_n310_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n674_), .A2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT114), .Z(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(new_n424_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n752_), .B2(new_n218_), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n747_), .B2(new_n634_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT115), .Z(new_n755_));
  NOR2_X1   g554(.A1(new_n578_), .A2(new_n219_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n751_), .B2(new_n756_), .ZN(G1337gat));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n641_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n641_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n758_), .A2(G99gat), .B1(new_n747_), .B2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g560(.A1(new_n747_), .A2(new_n227_), .A3(new_n651_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n750_), .A2(new_n651_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G106gat), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT52), .B(new_n227_), .C1(new_n750_), .C2(new_n651_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g567(.A1(new_n651_), .A2(new_n634_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n424_), .A3(new_n641_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n317_), .A2(new_n313_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT117), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n313_), .B1(new_n317_), .B2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n315_), .A2(KEYINPUT116), .A3(new_n316_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n777_), .A2(new_n778_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n322_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT121), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n323_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT56), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n784_), .A3(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n598_), .A2(new_n603_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n599_), .A2(KEYINPUT119), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n601_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n599_), .A2(KEYINPUT119), .ZN(new_n791_));
  OAI221_X1 g590(.A(new_n611_), .B1(new_n601_), .B2(new_n788_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n605_), .A2(new_n608_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n793_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n325_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n787_), .A2(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n781_), .A2(new_n784_), .A3(new_n782_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n771_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT58), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n771_), .B(new_n803_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n802_), .A2(new_n285_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n624_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n613_), .A2(new_n326_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n785_), .A2(KEYINPUT56), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(KEYINPUT118), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n783_), .A2(new_n810_), .A3(new_n786_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n797_), .B1(new_n328_), .B2(new_n326_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT57), .B(new_n806_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(new_n797_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n809_), .A2(new_n811_), .B1(new_n329_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n815_), .B1(new_n817_), .B2(new_n624_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n310_), .B1(new_n805_), .B2(new_n819_), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n335_), .A2(KEYINPUT54), .A3(new_n613_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT54), .B1(new_n335_), .B2(new_n613_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n770_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n613_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n718_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n826_), .B1(new_n829_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g629(.A(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n334_), .B2(KEYINPUT60), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n824_), .B(new_n832_), .C1(KEYINPUT60), .C2(new_n831_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n334_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n831_), .ZN(G1341gat));
  INV_X1    g634(.A(G127gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n824_), .A2(new_n836_), .A3(new_n309_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n310_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n836_), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n627_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n824_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n285_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n844_), .B2(new_n840_), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n651_), .A2(new_n375_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n578_), .A2(new_n424_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n814_), .A2(new_n818_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n802_), .A2(new_n285_), .A3(new_n804_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n309_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n823_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n847_), .B(new_n849_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n718_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n384_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n334_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n385_), .ZN(G1345gat));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT123), .B1(new_n854_), .B2(new_n310_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n854_), .A2(KEYINPUT123), .A3(new_n310_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n863_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n861_), .A3(new_n859_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(new_n854_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G162gat), .B1(new_n868_), .B2(new_n841_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n663_), .A2(new_n668_), .A3(G162gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(new_n870_), .ZN(G1347gat));
  NAND2_X1  g670(.A1(new_n820_), .A2(new_n823_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n578_), .A2(new_n424_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(new_n651_), .A3(new_n375_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(new_n613_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n876_), .A2(new_n877_), .A3(G169gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n872_), .A2(new_n875_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n534_), .A3(new_n613_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n876_), .B2(G169gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n878_), .B1(new_n881_), .B2(new_n882_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n879_), .A2(new_n334_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n518_), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n879_), .A2(new_n310_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n363_), .C1(KEYINPUT124), .C2(G183gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(G183gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n886_), .B2(new_n889_), .ZN(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n879_), .B2(new_n843_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n841_), .A2(new_n538_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n879_), .B2(new_n892_), .ZN(G1351gat));
  AOI211_X1 g692(.A(new_n846_), .B(new_n874_), .C1(new_n820_), .C2(new_n823_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n613_), .C1(KEYINPUT125), .C2(G197gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT125), .B(G197gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n872_), .A2(new_n847_), .A3(new_n873_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n718_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1352gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n334_), .ZN(new_n900_));
  AND2_X1   g699(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n902_), .ZN(G1353gat));
  AOI211_X1 g703(.A(KEYINPUT63), .B(G211gat), .C1(new_n894_), .C2(new_n309_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT63), .B(G211gat), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n897_), .A2(new_n310_), .A3(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1354gat));
  AOI21_X1  g707(.A(new_n441_), .B1(new_n894_), .B2(new_n285_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n627_), .A2(G218gat), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n897_), .A2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT127), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G218gat), .B1(new_n897_), .B2(new_n843_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n894_), .A2(new_n910_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n913_), .A2(new_n917_), .ZN(G1355gat));
endmodule


