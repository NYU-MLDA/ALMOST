//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n987_, new_n988_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1012_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1022_, new_n1023_, new_n1024_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT81), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n203_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n213_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n212_), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222_));
  OAI221_X1 g021(.A(new_n221_), .B1(G183gat), .B2(G190gat), .C1(new_n213_), .C2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n218_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n215_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n211_), .A2(new_n220_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT30), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n226_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n209_), .A2(new_n210_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT78), .B1(new_n207_), .B2(new_n208_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n220_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT30), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n228_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G71gat), .ZN(new_n240_));
  INV_X1    g039(.A(G99gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n228_), .A2(new_n235_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n206_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT80), .B(G43gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT31), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n243_), .A2(new_n245_), .A3(new_n206_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n249_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(new_n253_), .B2(new_n246_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G8gat), .B(G36gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(G64gat), .B(G92gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G226gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT19), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n226_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n221_), .B1(new_n213_), .B2(new_n222_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n217_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n207_), .A2(KEYINPUT93), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(G183gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT25), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n276_), .A3(new_n208_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT94), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n219_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n269_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n277_), .B2(new_n219_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n266_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT96), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G204gat), .ZN(new_n286_));
  INV_X1    g085(.A(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G197gat), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(new_n285_), .A3(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT21), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n289_), .B2(KEYINPUT90), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n286_), .A2(new_n288_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n290_), .B1(new_n298_), .B2(KEYINPUT21), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n293_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  OAI211_X1 g100(.A(KEYINPUT21), .B(new_n295_), .C1(new_n298_), .C2(new_n294_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT91), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n292_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n277_), .A2(new_n219_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT94), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n279_), .A3(new_n269_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(KEYINPUT96), .A3(new_n266_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n284_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT20), .ZN(new_n310_));
  INV_X1    g109(.A(new_n292_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT91), .B1(new_n301_), .B2(new_n302_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n297_), .A2(new_n293_), .A3(new_n299_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n314_), .B2(new_n233_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n264_), .B1(new_n309_), .B2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n304_), .B1(new_n307_), .B2(new_n266_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT20), .B1(new_n314_), .B2(new_n233_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n263_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n261_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n263_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n307_), .A2(new_n304_), .A3(new_n266_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n322_), .A3(new_n264_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n323_), .A3(new_n260_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(KEYINPUT27), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT27), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n321_), .A2(new_n323_), .A3(new_n260_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n260_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT87), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT85), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT84), .B1(new_n340_), .B2(KEYINPUT85), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n345_), .A2(KEYINPUT86), .A3(KEYINPUT2), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n348_), .A2(new_n349_), .B1(G141gat), .B2(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n335_), .B1(new_n344_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT83), .B1(new_n334_), .B2(KEYINPUT1), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n333_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n357_), .B2(new_n334_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n345_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(new_n337_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n334_), .B1(new_n332_), .B2(KEYINPUT1), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(KEYINPUT83), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n331_), .B1(new_n354_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n357_), .A2(new_n365_), .A3(new_n334_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n361_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n366_), .B(new_n360_), .C1(new_n367_), .C2(new_n355_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n341_), .A2(new_n343_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n368_), .B(KEYINPUT87), .C1(new_n369_), .C2(new_n335_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT89), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n364_), .A2(new_n370_), .A3(new_n374_), .A4(KEYINPUT29), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n304_), .B1(G228gat), .B2(G233gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n354_), .A2(new_n363_), .ZN(new_n378_));
  XOR2_X1   g177(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n379_));
  OAI21_X1  g178(.A(new_n314_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(G228gat), .A3(G233gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G78gat), .B(G106gat), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G22gat), .B(G50gat), .Z(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n371_), .A2(new_n372_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n390_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n385_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n388_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n383_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n377_), .A2(new_n381_), .A3(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n384_), .A2(new_n391_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n394_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n377_), .A2(new_n381_), .A3(new_n395_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n395_), .B1(new_n377_), .B2(new_n381_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n203_), .A2(new_n205_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n202_), .A2(KEYINPUT81), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n202_), .A2(KEYINPUT81), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n204_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n364_), .A2(new_n407_), .A3(new_n370_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n206_), .A2(new_n378_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  AND3_X1   g214(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT4), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n364_), .A2(new_n407_), .A3(new_n370_), .A4(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n410_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n411_), .B(new_n415_), .C1(new_n416_), .C2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT4), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n419_), .A3(new_n418_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n415_), .B1(new_n424_), .B2(new_n411_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  AND4_X1   g225(.A1(new_n255_), .A2(new_n330_), .A3(new_n402_), .A4(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n397_), .A2(new_n401_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n323_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n282_), .A2(new_n314_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n310_), .B1(new_n227_), .B2(new_n304_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n264_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n261_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT27), .B1(new_n433_), .B2(new_n324_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n411_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n415_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n421_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n428_), .A2(KEYINPUT97), .A3(new_n325_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n309_), .A2(new_n315_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n263_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n319_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n260_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n324_), .A2(KEYINPUT27), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n329_), .B(new_n426_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n441_), .B1(new_n447_), .B2(new_n402_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n321_), .A2(new_n323_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n435_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n424_), .A2(KEYINPUT33), .A3(new_n411_), .A4(new_n415_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n433_), .A3(new_n455_), .A4(new_n324_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n423_), .A2(new_n418_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n410_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n408_), .A2(new_n409_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n453_), .B1(new_n459_), .B2(new_n419_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n415_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  OAI22_X1  g260(.A1(new_n451_), .A2(new_n452_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n402_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n440_), .A2(new_n448_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n255_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT82), .B1(new_n251_), .B2(new_n254_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n427_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT77), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G36gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G29gat), .ZN(new_n475_));
  INV_X1    g274(.A(G29gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(G36gat), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n475_), .A2(new_n477_), .A3(KEYINPUT71), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT71), .B1(new_n475_), .B2(new_n477_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n473_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n477_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT71), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n477_), .A3(KEYINPUT71), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n472_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT74), .B(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(G22gat), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  INV_X1    g292(.A(G22gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G8gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n489_), .A2(new_n492_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n492_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT74), .B(G1gat), .Z(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n486_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n486_), .B1(new_n497_), .B2(new_n503_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n471_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n497_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n480_), .A2(new_n485_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(KEYINPUT77), .A3(new_n504_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n507_), .A2(new_n509_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n480_), .A2(new_n485_), .A3(KEYINPUT15), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(new_n510_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n508_), .A3(new_n512_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G169gat), .B(G197gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  AND3_X1   g322(.A1(new_n514_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n514_), .B2(new_n520_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n470_), .A2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(G230gat), .A2(G233gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT11), .ZN(new_n529_));
  INV_X1    g328(.A(G64gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(G57gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(G57gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(G71gat), .ZN(new_n536_));
  INV_X1    g335(.A(G71gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT65), .ZN(new_n538_));
  OAI21_X1  g337(.A(G78gat), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(G57gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G64gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n531_), .A2(new_n541_), .A3(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(KEYINPUT65), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n535_), .A2(G71gat), .ZN(new_n544_));
  INV_X1    g343(.A(G78gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n534_), .A2(new_n539_), .A3(new_n542_), .A4(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n532_), .A2(new_n533_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT11), .B(new_n548_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n554_));
  INV_X1    g353(.A(G106gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n241_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n556_), .A2(new_n559_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT8), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT64), .ZN(new_n564_));
  AND2_X1   g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(KEYINPUT64), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n572_));
  AND3_X1   g371(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n555_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(G85gat), .ZN(new_n579_));
  INV_X1    g378(.A(G92gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT9), .A3(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n582_), .A2(KEYINPUT9), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n575_), .A2(new_n578_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n571_), .A2(new_n572_), .A3(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT66), .B1(new_n553_), .B2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n562_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n588_));
  AND4_X1   g387(.A1(new_n575_), .A2(new_n578_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n569_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT66), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(new_n552_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n591_), .A2(new_n552_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n528_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n591_), .B2(new_n552_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n528_), .B1(new_n591_), .B2(new_n552_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n547_), .A2(new_n551_), .A3(KEYINPUT68), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT68), .B1(new_n547_), .B2(new_n551_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT12), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT67), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n571_), .A2(KEYINPUT67), .A3(new_n572_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n589_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n598_), .B(new_n599_), .C1(new_n602_), .C2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n596_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT5), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT69), .Z(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n596_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT13), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT13), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n617_), .A2(KEYINPUT70), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT70), .B1(new_n617_), .B2(new_n618_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT34), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT72), .B1(new_n586_), .B2(new_n486_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n588_), .A2(new_n590_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT72), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n511_), .A4(new_n585_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n606_), .A2(new_n518_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT35), .B(new_n624_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G190gat), .B(G218gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(KEYINPUT36), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n604_), .A2(new_n605_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n585_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n517_), .A3(new_n516_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n631_), .A2(new_n635_), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n634_), .B(KEYINPUT36), .Z(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n631_), .B2(new_n642_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n643_), .A2(new_n646_), .A3(KEYINPUT37), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n638_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n641_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n644_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n631_), .A2(new_n635_), .A3(new_n642_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n647_), .A2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT76), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G127gat), .B(G155gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G183gat), .B(G211gat), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n658_), .B(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT17), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n658_), .B(new_n659_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT17), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n510_), .B(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(new_n553_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n553_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n662_), .A2(new_n665_), .A3(new_n668_), .A4(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n600_), .A2(new_n601_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n667_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(new_n671_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n672_), .A2(KEYINPUT17), .A3(new_n661_), .A4(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n670_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n654_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n622_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n527_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT38), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n438_), .A2(new_n487_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT98), .B1(new_n643_), .B2(new_n646_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n651_), .A2(new_n683_), .A3(new_n652_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n470_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n675_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n622_), .A2(new_n526_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G1gat), .B1(new_n690_), .B2(new_n426_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n679_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n681_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT99), .ZN(G1324gat));
  NAND2_X1  g493(.A1(new_n325_), .A2(new_n329_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n695_), .A3(new_n689_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G8gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT100), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(new_n699_), .A3(G8gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n700_), .A3(KEYINPUT39), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n678_), .A2(G8gat), .A3(new_n330_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT39), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n699_), .B1(new_n696_), .B2(G8gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n701_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1325gat));
  INV_X1    g508(.A(new_n678_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n238_), .A3(new_n468_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G15gat), .B1(new_n690_), .B2(new_n469_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n713_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(G1326gat));
  NAND3_X1  g515(.A1(new_n710_), .A2(new_n494_), .A3(new_n428_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G22gat), .B1(new_n690_), .B2(new_n402_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n718_), .A2(KEYINPUT103), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(KEYINPUT103), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n721_));
  AND3_X1   g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n717_), .B1(new_n722_), .B2(new_n723_), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n686_), .A2(new_n688_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n622_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n527_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G29gat), .B1(new_n728_), .B2(new_n438_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n526_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n621_), .A2(new_n730_), .A3(new_n688_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n470_), .B2(new_n654_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n647_), .A2(new_n653_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n439_), .A2(new_n397_), .A3(new_n401_), .A4(new_n325_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n735_), .A2(new_n441_), .B1(new_n462_), .B2(new_n402_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n468_), .B1(new_n736_), .B2(new_n440_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n733_), .B(new_n734_), .C1(new_n737_), .C2(new_n427_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n731_), .B1(new_n732_), .B2(new_n738_), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n476_), .B(new_n426_), .C1(new_n739_), .C2(KEYINPUT44), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n739_), .A2(KEYINPUT44), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n729_), .B1(new_n740_), .B2(new_n741_), .ZN(G1328gat));
  NAND2_X1  g541(.A1(new_n739_), .A2(KEYINPUT44), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n695_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n739_), .A2(KEYINPUT44), .ZN(new_n745_));
  OAI21_X1  g544(.A(G36gat), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n330_), .A2(G36gat), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n727_), .A2(KEYINPUT45), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT45), .B1(new_n727_), .B2(new_n748_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n746_), .A2(KEYINPUT46), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n330_), .B1(new_n739_), .B2(KEYINPUT44), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n474_), .B1(new_n741_), .B2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n749_), .A2(new_n750_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n752_), .A2(new_n757_), .ZN(G1329gat));
  INV_X1    g557(.A(G43gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n727_), .B2(new_n469_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n743_), .A2(G43gat), .A3(new_n255_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n745_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT47), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n760_), .C1(new_n761_), .C2(new_n745_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1330gat));
  AOI21_X1  g565(.A(G50gat), .B1(new_n728_), .B2(new_n428_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n743_), .A2(G50gat), .A3(new_n428_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n741_), .ZN(G1331gat));
  NAND2_X1  g568(.A1(new_n675_), .A2(new_n526_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n621_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n687_), .A2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(new_n540_), .A3(new_n426_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n464_), .A2(new_n469_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n427_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n526_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n621_), .A2(new_n676_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(KEYINPUT104), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n778_), .A2(KEYINPUT104), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n777_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT105), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n438_), .B1(new_n781_), .B2(KEYINPUT105), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n540_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT106), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT106), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n786_), .B(new_n540_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n773_), .B1(new_n785_), .B2(new_n787_), .ZN(G1332gat));
  NAND3_X1  g587(.A1(new_n781_), .A2(new_n530_), .A3(new_n695_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G64gat), .B1(new_n772_), .B2(new_n330_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(KEYINPUT48), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(KEYINPUT48), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(G1333gat));
  NAND3_X1  g592(.A1(new_n781_), .A2(new_n537_), .A3(new_n468_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G71gat), .B1(new_n772_), .B2(new_n469_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(KEYINPUT49), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(KEYINPUT49), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n796_), .B2(new_n797_), .ZN(G1334gat));
  NAND3_X1  g597(.A1(new_n781_), .A2(new_n545_), .A3(new_n428_), .ZN(new_n799_));
  OAI21_X1  g598(.A(G78gat), .B1(new_n772_), .B2(new_n402_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(KEYINPUT50), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(KEYINPUT50), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n799_), .B1(new_n801_), .B2(new_n802_), .ZN(G1335gat));
  NOR2_X1   g602(.A1(new_n470_), .A2(new_n730_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n621_), .A2(new_n725_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n438_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n621_), .A2(new_n730_), .A3(new_n675_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n732_), .B2(new_n738_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n426_), .A2(new_n579_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT108), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n810_), .A2(new_n579_), .B1(new_n813_), .B2(new_n815_), .ZN(G1336gat));
  OAI211_X1 g615(.A(new_n580_), .B(new_n695_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n813_), .A2(new_n695_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n580_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1337gat));
  NAND3_X1  g620(.A1(new_n255_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n809_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n807_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n241_), .B1(new_n813_), .B2(new_n468_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n826_), .B(new_n828_), .ZN(G1338gat));
  OAI211_X1 g628(.A(new_n555_), .B(new_n428_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n830_));
  AOI211_X1 g629(.A(KEYINPUT52), .B(new_n555_), .C1(new_n813_), .C2(new_n428_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n733_), .B1(new_n776_), .B2(new_n734_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n470_), .A2(KEYINPUT43), .A3(new_n654_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n428_), .B(new_n811_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n835_), .B2(G106gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n830_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT53), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n830_), .B(new_n839_), .C1(new_n831_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1339gat));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n770_), .B1(new_n618_), .B2(new_n617_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n654_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n843_), .B2(new_n654_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(KEYINPUT111), .A2(KEYINPUT58), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n598_), .B1(new_n602_), .B2(new_n606_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n528_), .B1(new_n849_), .B2(new_n594_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT68), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n552_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n547_), .A2(new_n551_), .A3(KEYINPUT68), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n597_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n637_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n855_), .A2(KEYINPUT55), .A3(new_n598_), .A4(new_n599_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n607_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n850_), .A2(new_n856_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n613_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(KEYINPUT56), .A3(new_n613_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n514_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n507_), .A2(new_n508_), .A3(new_n513_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n506_), .A2(new_n508_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n523_), .B1(new_n519_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n615_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n848_), .B1(new_n864_), .B2(new_n872_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n859_), .A2(KEYINPUT56), .A3(new_n613_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n859_), .B2(new_n613_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n872_), .B(new_n848_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n734_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT112), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n848_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n654_), .B1(new_n882_), .B2(new_n876_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n615_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n870_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n685_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n685_), .B(KEYINPUT57), .C1(new_n887_), .C2(new_n888_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n879_), .A2(new_n885_), .A3(new_n891_), .A4(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n847_), .B1(new_n893_), .B2(new_n688_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n428_), .A2(new_n695_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n255_), .A3(new_n438_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n842_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n891_), .B(new_n892_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n878_), .A2(KEYINPUT112), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n688_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n847_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n896_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(KEYINPUT113), .A3(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n897_), .A2(new_n904_), .A3(new_n730_), .ZN(new_n905_));
  INV_X1    g704(.A(G113gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT114), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n905_), .A2(KEYINPUT114), .A3(new_n906_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT59), .B1(new_n894_), .B2(new_n896_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n903_), .A2(KEYINPUT115), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n903_), .A2(KEYINPUT115), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n912_), .A2(new_n913_), .A3(KEYINPUT59), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n878_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n901_), .B1(new_n675_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n911_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT116), .B(G113gat), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n526_), .A2(new_n920_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n909_), .A2(new_n910_), .B1(new_n919_), .B2(new_n921_), .ZN(G1340gat));
  AND2_X1   g721(.A1(new_n897_), .A2(new_n904_), .ZN(new_n923_));
  INV_X1    g722(.A(G120gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n621_), .B2(KEYINPUT60), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n923_), .B(new_n925_), .C1(KEYINPUT60), .C2(new_n924_), .ZN(new_n926_));
  OAI21_X1  g725(.A(KEYINPUT117), .B1(new_n918_), .B2(new_n621_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(G120gat), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n918_), .A2(KEYINPUT117), .A3(new_n621_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n926_), .B1(new_n928_), .B2(new_n929_), .ZN(G1341gat));
  NAND3_X1  g729(.A1(new_n897_), .A2(new_n904_), .A3(new_n675_), .ZN(new_n931_));
  INV_X1    g730(.A(G127gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n911_), .A2(G127gat), .A3(new_n675_), .A4(new_n917_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n933_), .A2(KEYINPUT118), .A3(new_n934_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1342gat));
  INV_X1    g738(.A(G134gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n923_), .A2(new_n940_), .A3(new_n686_), .ZN(new_n941_));
  OAI21_X1  g740(.A(G134gat), .B1(new_n918_), .B2(new_n654_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1343gat));
  NAND2_X1  g742(.A1(new_n469_), .A2(new_n428_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n944_), .A2(new_n426_), .A3(new_n695_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n902_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n526_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(KEYINPUT119), .B(G141gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1344gat));
  INV_X1    g748(.A(new_n946_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n622_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g751(.A1(new_n946_), .A2(new_n688_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT61), .B(G155gat), .Z(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1346gat));
  AOI21_X1  g754(.A(G162gat), .B1(new_n950_), .B2(new_n686_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n734_), .A2(G162gat), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT120), .Z(new_n958_));
  AOI21_X1  g757(.A(new_n956_), .B1(new_n950_), .B2(new_n958_), .ZN(G1347gat));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n330_), .A2(new_n438_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n469_), .A2(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n916_), .A2(new_n402_), .A3(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n526_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n960_), .B1(new_n965_), .B2(new_n214_), .ZN(new_n966_));
  OAI211_X1 g765(.A(KEYINPUT62), .B(G169gat), .C1(new_n964_), .C2(new_n526_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n225_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n966_), .A2(new_n967_), .A3(new_n968_), .ZN(G1348gat));
  INV_X1    g768(.A(new_n964_), .ZN(new_n970_));
  AOI21_X1  g769(.A(G176gat), .B1(new_n970_), .B2(new_n622_), .ZN(new_n971_));
  OAI21_X1  g770(.A(KEYINPUT121), .B1(new_n894_), .B2(new_n428_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n902_), .A2(new_n973_), .A3(new_n402_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n972_), .A2(new_n974_), .ZN(new_n975_));
  NOR4_X1   g774(.A1(new_n621_), .A2(new_n469_), .A3(new_n962_), .A4(new_n215_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n971_), .B1(new_n975_), .B2(new_n976_), .ZN(G1349gat));
  NAND2_X1  g776(.A1(new_n270_), .A2(new_n276_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n970_), .A2(new_n978_), .A3(new_n675_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n963_), .A2(new_n675_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n980_), .B1(new_n972_), .B2(new_n974_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n979_), .B1(new_n981_), .B2(G183gat), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(KEYINPUT122), .ZN(new_n983_));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n984_));
  OAI211_X1 g783(.A(new_n979_), .B(new_n984_), .C1(new_n981_), .C2(G183gat), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n983_), .A2(new_n985_), .ZN(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n964_), .B2(new_n654_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n686_), .A2(new_n208_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n987_), .B1(new_n964_), .B2(new_n988_), .ZN(G1351gat));
  NOR2_X1   g788(.A1(new_n944_), .A2(new_n962_), .ZN(new_n990_));
  INV_X1    g789(.A(new_n990_), .ZN(new_n991_));
  NOR3_X1   g790(.A1(new_n894_), .A2(new_n526_), .A3(new_n991_), .ZN(new_n992_));
  OAI21_X1  g791(.A(KEYINPUT124), .B1(new_n992_), .B2(G197gat), .ZN(new_n993_));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n902_), .A2(new_n990_), .ZN(new_n995_));
  OAI211_X1 g794(.A(new_n994_), .B(new_n285_), .C1(new_n995_), .C2(new_n526_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n993_), .A2(new_n996_), .ZN(new_n997_));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n998_));
  NOR2_X1   g797(.A1(new_n894_), .A2(new_n991_), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n526_), .A2(new_n285_), .ZN(new_n1000_));
  AOI21_X1  g799(.A(new_n998_), .B1(new_n999_), .B2(new_n1000_), .ZN(new_n1001_));
  INV_X1    g800(.A(new_n1000_), .ZN(new_n1002_));
  NOR4_X1   g801(.A1(new_n894_), .A2(KEYINPUT123), .A3(new_n991_), .A4(new_n1002_), .ZN(new_n1003_));
  NOR2_X1   g802(.A1(new_n1001_), .A2(new_n1003_), .ZN(new_n1004_));
  OAI21_X1  g803(.A(KEYINPUT125), .B1(new_n997_), .B2(new_n1004_), .ZN(new_n1005_));
  INV_X1    g804(.A(new_n1003_), .ZN(new_n1006_));
  OAI21_X1  g805(.A(KEYINPUT123), .B1(new_n995_), .B2(new_n1002_), .ZN(new_n1007_));
  NAND2_X1  g806(.A1(new_n1006_), .A2(new_n1007_), .ZN(new_n1008_));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n1009_));
  NAND4_X1  g808(.A1(new_n1008_), .A2(new_n1009_), .A3(new_n993_), .A4(new_n996_), .ZN(new_n1010_));
  NAND2_X1  g809(.A1(new_n1005_), .A2(new_n1010_), .ZN(G1352gat));
  NAND2_X1  g810(.A1(new_n999_), .A2(new_n622_), .ZN(new_n1012_));
  XNOR2_X1  g811(.A(new_n1012_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g812(.A(new_n688_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1014_));
  INV_X1    g813(.A(new_n1014_), .ZN(new_n1015_));
  OAI21_X1  g814(.A(KEYINPUT126), .B1(new_n995_), .B2(new_n1015_), .ZN(new_n1016_));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1017_));
  NAND3_X1  g816(.A1(new_n999_), .A2(new_n1017_), .A3(new_n1014_), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(new_n1016_), .A2(new_n1018_), .ZN(new_n1019_));
  NOR2_X1   g818(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1020_));
  XOR2_X1   g819(.A(new_n1019_), .B(new_n1020_), .Z(G1354gat));
  XOR2_X1   g820(.A(KEYINPUT127), .B(G218gat), .Z(new_n1022_));
  NOR3_X1   g821(.A1(new_n995_), .A2(new_n654_), .A3(new_n1022_), .ZN(new_n1023_));
  NAND2_X1  g822(.A1(new_n999_), .A2(new_n686_), .ZN(new_n1024_));
  AOI21_X1  g823(.A(new_n1023_), .B1(new_n1024_), .B2(new_n1022_), .ZN(G1355gat));
endmodule


