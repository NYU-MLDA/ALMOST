//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  AND4_X1   g010(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT8), .B1(new_n207_), .B2(new_n213_), .ZN(new_n214_));
  OR3_X1    g013(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n203_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n207_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n212_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G71gat), .B(G78gat), .Z(new_n222_));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n222_), .B1(KEYINPUT11), .B2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n224_), .A2(KEYINPUT67), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT67), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(KEYINPUT11), .A3(new_n223_), .A4(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n221_), .B(new_n231_), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT12), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT12), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n221_), .A2(new_n234_), .A3(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G230gat), .A2(G233gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT64), .Z(new_n238_));
  AND2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n232_), .A2(new_n238_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G120gat), .B(G148gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT5), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G176gat), .B(G204gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n241_), .A2(new_n245_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT13), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(KEYINPUT13), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G134gat), .B(G162gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(G190gat), .B(G218gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT36), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G29gat), .B(G36gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT69), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G43gat), .B(G50gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n221_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT71), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n220_), .B(new_n263_), .C1(new_n214_), .C2(new_n219_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G232gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT34), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT35), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(KEYINPUT73), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(KEYINPUT73), .B2(new_n274_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n267_), .A2(new_n268_), .A3(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT74), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n267_), .A2(new_n268_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n274_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT72), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n258_), .B(new_n259_), .C1(new_n279_), .C2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n285_), .A2(new_n257_), .A3(new_n256_), .A4(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT37), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(KEYINPUT37), .A3(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G1gat), .ZN(new_n292_));
  INV_X1    g091(.A(G8gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G1gat), .B(G8gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(new_n231_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G127gat), .B(G155gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G183gat), .B(G211gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT17), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  OR3_X1    g111(.A1(new_n304_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(KEYINPUT77), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT77), .B1(new_n304_), .B2(new_n311_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n291_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n253_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT78), .ZN(new_n321_));
  XOR2_X1   g120(.A(G1gat), .B(G29gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(G57gat), .B(G85gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G134gat), .Z(new_n328_));
  INV_X1    g127(.A(KEYINPUT84), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT84), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  INV_X1    g139(.A(G141gat), .ZN(new_n341_));
  INV_X1    g140(.A(G148gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT87), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT87), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n345_), .A2(new_n340_), .A3(new_n341_), .A4(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(KEYINPUT2), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT88), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n348_), .B(new_n349_), .C1(new_n351_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n347_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(KEYINPUT88), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n350_), .A2(KEYINPUT2), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n358_), .B1(new_n362_), .B2(new_n348_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n339_), .B1(new_n355_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n337_), .A2(new_n365_), .A3(new_n338_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n341_), .A2(new_n342_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n349_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT86), .B1(new_n367_), .B2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n368_), .A2(new_n349_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n366_), .A3(new_n373_), .A4(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT100), .B(KEYINPUT4), .Z(new_n377_));
  NAND3_X1  g176(.A1(new_n336_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n364_), .A2(new_n375_), .A3(KEYINPUT99), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT98), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n334_), .A2(new_n335_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT88), .B(KEYINPUT2), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT89), .B1(new_n386_), .B2(new_n359_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n387_), .A2(new_n347_), .A3(new_n358_), .A4(new_n354_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n388_), .A2(new_n339_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT98), .B1(new_n389_), .B2(KEYINPUT99), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n364_), .A2(new_n375_), .A3(KEYINPUT98), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n336_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n385_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n381_), .B1(new_n393_), .B2(KEYINPUT4), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n382_), .A2(new_n383_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n336_), .A3(new_n391_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n380_), .B1(new_n396_), .B2(new_n385_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n327_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n379_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n396_), .B2(new_n385_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n399_), .B(new_n326_), .C1(new_n401_), .C2(new_n381_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n376_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT28), .B1(new_n376_), .B2(KEYINPUT29), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G22gat), .B(G50gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G197gat), .B(G204gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT21), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G218gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G211gat), .ZN(new_n414_));
  INV_X1    g213(.A(G211gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G218gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n416_), .A3(KEYINPUT91), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n415_), .A2(G218gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n413_), .A2(G211gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n412_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n417_), .ZN(new_n423_));
  INV_X1    g222(.A(G197gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(G204gat), .ZN(new_n426_));
  INV_X1    g225(.A(G204gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G197gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT21), .B(new_n425_), .C1(new_n429_), .C2(KEYINPUT90), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n410_), .A2(new_n411_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n423_), .A2(new_n430_), .A3(KEYINPUT92), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n421_), .A2(new_n417_), .B1(new_n411_), .B2(new_n410_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT92), .B1(new_n434_), .B2(new_n430_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n422_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT93), .ZN(new_n437_));
  INV_X1    g236(.A(new_n422_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT92), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n414_), .A2(new_n416_), .A3(KEYINPUT91), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT91), .B1(new_n414_), .B2(new_n416_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n431_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n425_), .A2(KEYINPUT21), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT90), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n410_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n439_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n438_), .B1(new_n446_), .B2(new_n432_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT93), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n376_), .A2(KEYINPUT29), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n437_), .A2(new_n449_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n436_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(G228gat), .A3(G233gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G78gat), .B(G106gat), .Z(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n455_), .A2(new_n456_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n409_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n457_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n455_), .A2(new_n456_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n408_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G183gat), .A2(G190gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n467_));
  INV_X1    g266(.A(G169gat), .ZN(new_n468_));
  INV_X1    g267(.A(G176gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n466_), .B(new_n467_), .C1(new_n470_), .C2(KEYINPUT24), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(G169gat), .B2(G176gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT25), .B(G183gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476_));
  INV_X1    g275(.A(G190gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(KEYINPUT26), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT26), .B(G190gat), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n475_), .B(new_n478_), .C1(new_n479_), .C2(new_n476_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n466_), .B(new_n467_), .C1(G183gat), .C2(G190gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(new_n468_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n474_), .A2(new_n480_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486_));
  INV_X1    g285(.A(G43gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n485_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G227gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G15gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT30), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n384_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n491_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(new_n403_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G8gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT18), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G226gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n437_), .A2(new_n449_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(new_n485_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n471_), .B(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n473_), .B1(new_n479_), .B2(new_n475_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n483_), .B1(new_n481_), .B2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n481_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT97), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n436_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n512_), .A2(new_n513_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT97), .B1(new_n447_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n507_), .B1(new_n510_), .B2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n508_), .B1(new_n447_), .B2(new_n522_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n507_), .B(new_n526_), .C1(new_n509_), .C2(new_n485_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n503_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n446_), .A2(new_n432_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n448_), .B1(new_n530_), .B2(new_n422_), .ZN(new_n531_));
  AOI211_X1 g330(.A(KEYINPUT93), .B(new_n438_), .C1(new_n446_), .C2(new_n432_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n485_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n533_), .A3(KEYINPUT20), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n506_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(new_n527_), .A3(new_n502_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT27), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n531_), .A2(new_n532_), .A3(new_n485_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n526_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n506_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n524_), .A2(new_n533_), .A3(KEYINPUT20), .A4(new_n507_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n503_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n536_), .A3(KEYINPUT27), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT106), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n463_), .B(new_n498_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n403_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n539_), .A2(new_n552_), .A3(new_n546_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n502_), .A2(KEYINPUT32), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n544_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n535_), .A2(new_n527_), .A3(new_n554_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n403_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT103), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n403_), .A2(new_n556_), .A3(new_n557_), .A4(KEYINPUT103), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n393_), .A2(KEYINPUT4), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n378_), .A2(new_n379_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n326_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT102), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n393_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n396_), .A2(KEYINPUT102), .A3(new_n385_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n380_), .A3(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n402_), .A2(new_n562_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n394_), .A2(new_n397_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(KEYINPUT33), .A3(new_n326_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n570_), .A2(new_n529_), .A3(new_n536_), .A4(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n560_), .A2(new_n561_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n463_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT104), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n553_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(KEYINPUT104), .A3(new_n463_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n496_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT105), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n551_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n574_), .A2(KEYINPUT104), .A3(new_n463_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT104), .B1(new_n574_), .B2(new_n463_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n553_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n584_), .A2(KEYINPUT105), .A3(new_n496_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT79), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n263_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n301_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT80), .ZN(new_n590_));
  INV_X1    g389(.A(new_n301_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n265_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n588_), .A2(new_n301_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n597_), .B2(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT81), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n603_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT82), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n586_), .A2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n321_), .A2(new_n292_), .A3(new_n403_), .A4(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT107), .Z(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT38), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n283_), .A2(KEYINPUT108), .A3(new_n286_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT108), .B1(new_n283_), .B2(new_n286_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n586_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n251_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n615_), .A2(new_n606_), .A3(new_n317_), .A4(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n403_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n610_), .A2(KEYINPUT38), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n611_), .A2(new_n619_), .A3(new_n620_), .ZN(G1324gat));
  AOI21_X1  g420(.A(new_n293_), .B1(KEYINPUT109), .B2(KEYINPUT39), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n549_), .A2(new_n550_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n622_), .B1(new_n617_), .B2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(KEYINPUT109), .A2(KEYINPUT39), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  NAND2_X1  g426(.A1(new_n321_), .A2(new_n608_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n293_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n617_), .B2(new_n497_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT41), .Z(new_n633_));
  OR2_X1    g432(.A1(new_n497_), .A2(G15gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n628_), .B2(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n617_), .B2(new_n463_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n463_), .A2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n628_), .B2(new_n639_), .ZN(G1327gat));
  INV_X1    g439(.A(new_n614_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(new_n317_), .A3(new_n251_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n608_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT113), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n403_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT112), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  INV_X1    g446(.A(new_n606_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n251_), .A2(new_n648_), .A3(new_n317_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n291_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n653_), .B(new_n291_), .C1(new_n581_), .C2(new_n585_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n650_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT111), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n647_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT111), .B(new_n650_), .C1(new_n652_), .C2(new_n654_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n646_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n654_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT105), .B1(new_n584_), .B2(new_n496_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n577_), .A2(new_n578_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n580_), .A3(new_n497_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n663_), .A3(new_n551_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n653_), .B1(new_n664_), .B2(new_n291_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n649_), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT44), .B1(new_n666_), .B2(KEYINPUT111), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n655_), .A2(new_n656_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(KEYINPUT112), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n659_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n655_), .A2(KEYINPUT44), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n403_), .A2(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n645_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n644_), .A2(new_n675_), .A3(new_n623_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT114), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n671_), .A2(new_n623_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n657_), .A2(new_n646_), .A3(new_n658_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT112), .B1(new_n667_), .B2(new_n668_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n678_), .B(new_n680_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G36gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n679_), .B1(new_n659_), .B2(new_n669_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n678_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n677_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT115), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(KEYINPUT115), .A2(KEYINPUT46), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n687_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n670_), .A2(new_n680_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT114), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n675_), .B1(new_n685_), .B2(new_n678_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n696_), .A2(new_n688_), .A3(new_n689_), .A4(new_n677_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n692_), .A2(new_n697_), .ZN(G1329gat));
  AOI21_X1  g497(.A(G43gat), .B1(new_n644_), .B2(new_n496_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n497_), .A2(new_n487_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n672_), .B2(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g501(.A(new_n463_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G50gat), .B1(new_n644_), .B2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(G50gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n672_), .B2(new_n705_), .ZN(G1331gat));
  INV_X1    g505(.A(new_n253_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n707_), .A2(new_n607_), .A3(new_n317_), .A4(new_n615_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n618_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n586_), .A2(new_n606_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n319_), .A3(new_n251_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n618_), .A2(G57gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT116), .Z(G1332gat));
  OAI21_X1  g513(.A(G64gat), .B1(new_n708_), .B2(new_n624_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT48), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n624_), .A2(G64gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n711_), .B2(new_n717_), .ZN(G1333gat));
  OAI21_X1  g517(.A(G71gat), .B1(new_n708_), .B2(new_n497_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT49), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n497_), .A2(G71gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT117), .Z(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n711_), .B2(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n708_), .B2(new_n463_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n463_), .A2(G78gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n711_), .B2(new_n726_), .ZN(G1335gat));
  NOR3_X1   g526(.A1(new_n253_), .A2(new_n317_), .A3(new_n641_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n710_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n209_), .A3(new_n403_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n251_), .A2(new_n648_), .A3(new_n318_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT118), .Z(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n403_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n735_), .B2(new_n209_), .ZN(G1336gat));
  OAI21_X1  g535(.A(new_n210_), .B1(new_n729_), .B2(new_n624_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT119), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n624_), .A2(new_n210_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n734_), .B2(new_n739_), .ZN(G1337gat));
  NAND2_X1  g539(.A1(new_n734_), .A2(new_n496_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n496_), .A2(new_n204_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n741_), .A2(G99gat), .B1(new_n730_), .B2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g543(.A(new_n205_), .B1(new_n734_), .B2(new_n703_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT52), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n730_), .A2(new_n205_), .A3(new_n703_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g548(.A1(new_n648_), .A2(new_n246_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n245_), .B1(new_n239_), .B2(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n239_), .A2(new_n751_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n236_), .A2(new_n238_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n597_), .A2(new_n594_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n593_), .A2(new_n594_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n602_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n602_), .B2(new_n598_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n248_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n641_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(KEYINPUT57), .A3(new_n641_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n291_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n762_), .A2(new_n246_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n757_), .A2(new_n769_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT58), .Z(new_n771_));
  OAI211_X1 g570(.A(new_n766_), .B(new_n767_), .C1(new_n768_), .C2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n318_), .ZN(new_n773_));
  AND4_X1   g572(.A1(new_n607_), .A2(new_n317_), .A3(new_n250_), .A4(new_n249_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n768_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(KEYINPUT120), .A2(KEYINPUT54), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT120), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n774_), .B(new_n768_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(KEYINPUT121), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT121), .B1(new_n780_), .B2(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n773_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n623_), .A2(new_n497_), .A3(new_n703_), .A4(new_n618_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G113gat), .B1(new_n786_), .B2(new_n606_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n784_), .A2(KEYINPUT59), .A3(new_n785_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT59), .B1(new_n784_), .B2(new_n785_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT122), .B(G113gat), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n607_), .A2(new_n792_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT123), .Z(new_n794_));
  AOI21_X1  g593(.A(new_n787_), .B1(new_n791_), .B2(new_n794_), .ZN(G1340gat));
  XNOR2_X1  g594(.A(KEYINPUT124), .B(G120gat), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n251_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n784_), .B(new_n785_), .C1(KEYINPUT60), .C2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n798_), .B2(KEYINPUT60), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n707_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n790_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT125), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT125), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n799_), .B(new_n803_), .C1(new_n790_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1341gat));
  OAI21_X1  g604(.A(G127gat), .B1(new_n790_), .B2(new_n318_), .ZN(new_n806_));
  INV_X1    g605(.A(G127gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n786_), .A2(new_n807_), .A3(new_n317_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1342gat));
  AOI21_X1  g608(.A(G134gat), .B1(new_n786_), .B2(new_n614_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n291_), .A2(G134gat), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(KEYINPUT126), .Z(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n791_), .B2(new_n812_), .ZN(G1343gat));
  NOR3_X1   g612(.A1(new_n623_), .A2(new_n463_), .A3(new_n618_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n784_), .A2(new_n497_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n606_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n707_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g618(.A(KEYINPUT61), .B(G155gat), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT127), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n815_), .A2(new_n822_), .A3(new_n317_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n815_), .B2(new_n317_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n825_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n823_), .A3(new_n820_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1346gat));
  INV_X1    g628(.A(new_n815_), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n830_), .A2(G162gat), .A3(new_n641_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G162gat), .B1(new_n830_), .B2(new_n768_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1347gat));
  AND3_X1   g632(.A1(new_n623_), .A2(new_n463_), .A3(new_n498_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n784_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n606_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT62), .B1(new_n837_), .B2(KEYINPUT22), .ZN(new_n838_));
  OAI21_X1  g637(.A(G169gat), .B1(new_n837_), .B2(KEYINPUT62), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n468_), .B2(new_n838_), .ZN(G1348gat));
  OAI21_X1  g640(.A(G176gat), .B1(new_n835_), .B2(new_n253_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n251_), .A2(new_n469_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n835_), .B2(new_n843_), .ZN(G1349gat));
  NOR2_X1   g643(.A1(new_n835_), .A2(new_n318_), .ZN(new_n845_));
  MUX2_X1   g644(.A(G183gat), .B(new_n475_), .S(new_n845_), .Z(G1350gat));
  OAI21_X1  g645(.A(G190gat), .B1(new_n835_), .B2(new_n768_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n614_), .A2(new_n479_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n835_), .B2(new_n848_), .ZN(G1351gat));
  NAND4_X1  g648(.A1(new_n784_), .A2(new_n497_), .A3(new_n552_), .A4(new_n623_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n648_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n424_), .ZN(G1352gat));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n253_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n427_), .ZN(G1353gat));
  NOR2_X1   g653(.A1(new_n850_), .A2(new_n318_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n856_));
  AND2_X1   g655(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n855_), .B2(new_n856_), .ZN(G1354gat));
  OAI21_X1  g658(.A(G218gat), .B1(new_n850_), .B2(new_n768_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n614_), .A2(new_n413_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n850_), .B2(new_n861_), .ZN(G1355gat));
endmodule


