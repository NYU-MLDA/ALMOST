//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT8), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT66), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT7), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  AOI211_X1 g012(.A(G99gat), .B(G106gat), .C1(new_n206_), .C2(KEYINPUT7), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n208_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n202_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n213_), .B1(new_n216_), .B2(KEYINPUT9), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT10), .B(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT9), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G85gat), .A3(G92gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(new_n220_), .B2(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n219_), .A2(new_n224_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n207_), .A2(new_n203_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(new_n203_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT8), .B(new_n216_), .C1(new_n231_), .C2(new_n213_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n218_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G57gat), .B(G64gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT11), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(KEYINPUT11), .ZN(new_n236_));
  XOR2_X1   g035(.A(G71gat), .B(G78gat), .Z(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n233_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n240_), .A2(new_n218_), .A3(new_n228_), .A4(new_n232_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(KEYINPUT12), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n245_), .A3(new_n241_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT64), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n242_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n243_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n249_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT67), .B(G204gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT5), .B(G176gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G120gat), .B(G148gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n255_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n255_), .A2(new_n261_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n262_), .A2(KEYINPUT13), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT13), .B1(new_n264_), .B2(new_n262_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT102), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G225gat), .A2(G233gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  OR3_X1    g075(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n278_));
  INV_X1    g077(.A(G141gat), .ZN(new_n279_));
  INV_X1    g078(.A(G148gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT3), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT83), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n283_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n283_), .A2(KEYINPUT85), .A3(new_n289_), .A4(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT84), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n297_), .B(new_n291_), .C1(new_n288_), .C2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n288_), .A2(new_n298_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT84), .B1(new_n301_), .B2(new_n290_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n299_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n273_), .A2(new_n275_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n281_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n306_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n296_), .A2(new_n305_), .A3(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT81), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT81), .B1(new_n309_), .B2(new_n311_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n296_), .B2(new_n305_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT4), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n296_), .A2(new_n305_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n314_), .A2(new_n315_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n270_), .B1(new_n318_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT97), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n313_), .A2(new_n317_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(new_n270_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n296_), .A2(new_n305_), .A3(new_n312_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n321_), .A2(new_n270_), .A3(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(KEYINPUT97), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n324_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G57gat), .B(G85gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT100), .B1(new_n331_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n270_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n322_), .B1(new_n321_), .B2(new_n328_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n317_), .A2(KEYINPUT4), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n326_), .A2(new_n325_), .A3(new_n270_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n329_), .A2(KEYINPUT97), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .A4(new_n337_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT100), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n336_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n338_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT27), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G92gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT18), .B(G64gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(G197gat), .B(G204gat), .Z(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(KEYINPUT21), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(KEYINPUT21), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(KEYINPUT24), .A3(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT25), .B(G183gat), .Z(new_n366_));
  AND2_X1   g165(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT77), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(KEYINPUT23), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n375_));
  INV_X1    g174(.A(new_n372_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n365_), .B(new_n380_), .C1(new_n366_), .C2(new_n369_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n371_), .A2(new_n377_), .A3(new_n379_), .A4(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n383_));
  OAI21_X1  g182(.A(G169gat), .B1(new_n383_), .B2(G176gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G169gat), .ZN(new_n386_));
  INV_X1    g185(.A(G176gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n376_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n376_), .B2(new_n375_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  OAI221_X1 g191(.A(new_n384_), .B1(new_n385_), .B2(new_n388_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n361_), .A2(new_n382_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n377_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n388_), .B(new_n364_), .C1(new_n395_), .C2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT94), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n377_), .B1(G183gat), .B2(G190gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT94), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n388_), .A4(new_n364_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n363_), .A2(KEYINPUT24), .A3(new_n364_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT91), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT26), .ZN(new_n405_));
  INV_X1    g204(.A(G190gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n366_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n402_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT92), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n366_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT92), .B1(new_n415_), .B2(new_n402_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n391_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n414_), .A2(new_n416_), .A3(new_n417_), .A4(new_n379_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT93), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n410_), .A2(new_n411_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n365_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n391_), .B1(new_n422_), .B2(KEYINPUT92), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n412_), .A2(new_n413_), .B1(new_n378_), .B2(new_n362_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT93), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n401_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT20), .B(new_n394_), .C1(new_n426_), .C2(new_n361_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT19), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT90), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n397_), .A2(new_n400_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n418_), .A2(new_n419_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT93), .B1(new_n423_), .B2(new_n424_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n361_), .B(new_n431_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n429_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n382_), .A2(new_n393_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n361_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n434_), .A2(KEYINPUT95), .A3(new_n435_), .A4(new_n439_), .ZN(new_n443_));
  AOI221_X4 g242(.A(new_n356_), .B1(new_n427_), .B2(new_n430_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n443_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n427_), .A2(new_n430_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n355_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n351_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G78gat), .B(G106gat), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G228gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n296_), .B2(new_n305_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n454_), .B2(new_n361_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n454_), .A2(new_n452_), .A3(new_n361_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n450_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n319_), .A2(KEYINPUT29), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n451_), .A3(new_n438_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n455_), .A3(new_n449_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(KEYINPUT88), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n460_), .A2(new_n455_), .A3(new_n463_), .A4(new_n449_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G22gat), .B(G50gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n296_), .A2(new_n305_), .A3(new_n453_), .A4(new_n467_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n464_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n469_), .A2(KEYINPUT87), .A3(new_n470_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n462_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n458_), .A2(KEYINPUT89), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n478_), .B(new_n450_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n477_), .A2(new_n479_), .A3(new_n461_), .A4(new_n471_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n437_), .A2(new_n438_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT98), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(KEYINPUT20), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n418_), .A2(new_n396_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT99), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n418_), .A2(KEYINPUT99), .A3(new_n396_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n484_), .B1(new_n489_), .B2(new_n361_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n436_), .A2(KEYINPUT98), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n435_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n427_), .A2(new_n430_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n356_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n429_), .B1(new_n426_), .B2(new_n361_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT95), .B1(new_n495_), .B2(new_n439_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n443_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n355_), .B(new_n446_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(KEYINPUT27), .A3(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n350_), .A2(new_n448_), .A3(new_n481_), .A4(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n446_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n356_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n270_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n326_), .A2(new_n339_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n336_), .A3(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n502_), .A2(new_n498_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n345_), .B(KEYINPUT33), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n427_), .A2(new_n430_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n490_), .A2(new_n491_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n508_), .B(new_n509_), .C1(new_n510_), .C2(new_n435_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n442_), .A2(new_n443_), .B1(new_n430_), .B2(new_n427_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n506_), .A2(new_n507_), .B1(new_n349_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n500_), .B1(new_n514_), .B2(new_n481_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n320_), .B(KEYINPUT30), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(new_n437_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n437_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G71gat), .B(G99gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G227gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G43gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n522_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n517_), .A2(new_n518_), .A3(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n523_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n481_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n531_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT101), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT27), .B1(new_n502_), .B2(new_n498_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n494_), .A2(KEYINPUT27), .A3(new_n498_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n448_), .A2(KEYINPUT101), .A3(new_n499_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n534_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n515_), .A2(new_n532_), .B1(new_n540_), .B2(new_n350_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G8gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT73), .ZN(new_n543_));
  XOR2_X1   g342(.A(G15gat), .B(G22gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT72), .B(G1gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G8gat), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n546_), .B2(KEYINPUT14), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n543_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G29gat), .B(G36gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT15), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT75), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n548_), .A2(new_n552_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT75), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n558_), .A3(new_n553_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n556_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n557_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n548_), .A2(new_n552_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(KEYINPUT76), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT76), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n269_), .B1(new_n541_), .B2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n507_), .A2(new_n498_), .A3(new_n502_), .A4(new_n505_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n349_), .A2(new_n513_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n481_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n448_), .A2(new_n499_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n481_), .A2(new_n345_), .A3(new_n338_), .A4(new_n348_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n532_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n534_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n536_), .A2(new_n537_), .A3(new_n535_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT101), .B1(new_n448_), .B2(new_n499_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n584_), .B(new_n350_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n575_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(KEYINPUT102), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n268_), .B1(new_n576_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n553_), .A2(new_n233_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n596_));
  INV_X1    g395(.A(new_n552_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n592_), .B(new_n596_), .C1(new_n597_), .C2(new_n233_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601_));
  INV_X1    g400(.A(G162gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT69), .B(G134gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT36), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n605_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n600_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT70), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n600_), .A2(KEYINPUT70), .A3(new_n610_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n608_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT71), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT37), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(KEYINPUT37), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(new_n617_), .A3(KEYINPUT37), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(G211gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT16), .B(G183gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n240_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(new_n548_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n626_), .B1(new_n629_), .B2(KEYINPUT17), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(KEYINPUT17), .B2(new_n626_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(KEYINPUT74), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n622_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n591_), .A2(new_n634_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n635_), .A2(new_n350_), .A3(new_n545_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT38), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n615_), .B(KEYINPUT103), .Z(new_n639_));
  NOR2_X1   g438(.A1(new_n268_), .A2(new_n572_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n588_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n633_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n350_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n636_), .A2(new_n637_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(new_n644_), .A3(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n538_), .A2(new_n539_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n648_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n641_), .A2(KEYINPUT104), .A3(new_n642_), .A4(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(G8gat), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n649_), .A2(new_n654_), .A3(G8gat), .A4(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n635_), .A2(G8gat), .A3(new_n648_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(KEYINPUT40), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n643_), .B2(new_n532_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n635_), .A2(G15gat), .A3(new_n532_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  OAI21_X1  g465(.A(G22gat), .B1(new_n643_), .B2(new_n533_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT42), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n533_), .A2(G22gat), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT105), .Z(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n635_), .B2(new_n670_), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n642_), .A2(new_n616_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT102), .B1(new_n588_), .B2(new_n589_), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n269_), .B(new_n575_), .C1(new_n583_), .C2(new_n587_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n267_), .B(new_n672_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n675_), .A2(G29gat), .A3(new_n350_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n622_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n541_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n588_), .A2(new_n679_), .A3(new_n622_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n633_), .A3(new_n640_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(KEYINPUT44), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n681_), .A2(new_n633_), .A3(new_n640_), .A4(new_n684_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n349_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT107), .B1(new_n689_), .B2(G29gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n676_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  NOR2_X1   g491(.A1(new_n648_), .A2(G36gat), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT108), .B1(new_n675_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n591_), .A2(new_n697_), .A3(new_n672_), .A4(new_n693_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n695_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n695_), .B2(new_n698_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n648_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n701_));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n699_), .A2(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI221_X1 g504(.A(KEYINPUT46), .B1(new_n701_), .B2(new_n702_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  INV_X1    g506(.A(new_n675_), .ZN(new_n708_));
  INV_X1    g507(.A(G43gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n531_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n532_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n709_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1330gat));
  INV_X1    g513(.A(G50gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(new_n715_), .A3(new_n481_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n533_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n715_), .ZN(G1331gat));
  INV_X1    g517(.A(new_n572_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n267_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n541_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n634_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n349_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n633_), .B1(new_n574_), .B2(new_n573_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n588_), .A2(new_n639_), .A3(new_n268_), .A4(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n349_), .A2(G57gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1332gat));
  OAI21_X1  g529(.A(G64gat), .B1(new_n727_), .B2(new_n648_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT48), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n648_), .A2(G64gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n723_), .B2(new_n733_), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n727_), .B2(new_n532_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n532_), .A2(G71gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n723_), .B2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n727_), .B2(new_n533_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n533_), .A2(G78gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n723_), .B2(new_n742_), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n721_), .A2(new_n642_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n681_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n350_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n722_), .A2(new_n672_), .ZN(new_n747_));
  INV_X1    g546(.A(G85gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n349_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT110), .ZN(G1336gat));
  AOI21_X1  g550(.A(G92gat), .B1(new_n747_), .B2(new_n650_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n745_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n650_), .A2(G92gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n745_), .B2(new_n532_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n747_), .A2(new_n221_), .A3(new_n531_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g558(.A(new_n679_), .B1(new_n588_), .B2(new_n622_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT43), .B(new_n677_), .C1(new_n583_), .C2(new_n587_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n481_), .B(new_n744_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT111), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n681_), .A2(new_n764_), .A3(new_n481_), .A4(new_n744_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(G106gat), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n763_), .A2(new_n765_), .A3(new_n768_), .A4(G106gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n747_), .A2(new_n223_), .A3(new_n481_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n774_), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n251_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n244_), .A2(new_n249_), .A3(new_n246_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n249_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT55), .B1(new_n781_), .B2(KEYINPUT113), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n780_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n261_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT114), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n783_), .A2(KEYINPUT114), .A3(new_n785_), .A4(new_n261_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n787_), .A2(new_n719_), .A3(new_n264_), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT115), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n264_), .A2(new_n262_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n555_), .A2(new_n561_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n556_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n567_), .A3(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n569_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n572_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n264_), .A4(new_n788_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n790_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n616_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n264_), .A2(new_n795_), .A3(KEYINPUT116), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n569_), .A2(new_n794_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n263_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n784_), .A2(KEYINPUT56), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n783_), .A2(new_n785_), .A3(new_n261_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n808_), .A2(KEYINPUT58), .A3(new_n809_), .A4(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n622_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n800_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n803_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n633_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n726_), .A2(new_n620_), .A3(new_n267_), .A4(new_n621_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT54), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n820_), .A2(KEYINPUT112), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n819_), .A2(KEYINPUT54), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(KEYINPUT112), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n818_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT117), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n818_), .A2(new_n824_), .A3(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n540_), .A2(new_n349_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830_), .B2(new_n719_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n829_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT118), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n832_), .B2(new_n829_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n800_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT57), .B1(new_n800_), .B2(new_n616_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n622_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n642_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n817_), .A2(new_n843_), .A3(new_n633_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n824_), .A3(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n837_), .A2(new_n845_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n834_), .A2(KEYINPUT118), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n834_), .B2(new_n830_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n589_), .A2(G113gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n831_), .B1(new_n850_), .B2(new_n851_), .ZN(G1340gat));
  OAI21_X1  g651(.A(G120gat), .B1(new_n849_), .B2(new_n267_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  AOI21_X1  g653(.A(G120gat), .B1(new_n268_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT121), .B1(new_n854_), .B2(G120gat), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n830_), .B(new_n857_), .C1(new_n855_), .C2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n853_), .A2(new_n859_), .ZN(G1341gat));
  NAND2_X1  g659(.A1(new_n826_), .A2(new_n828_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n633_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G127gat), .B1(new_n862_), .B2(new_n829_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n642_), .A2(G127gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n850_), .B2(new_n864_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n677_), .A2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n848_), .B(new_n867_), .C1(new_n830_), .C2(new_n834_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n639_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n826_), .A2(new_n869_), .A3(new_n828_), .A4(new_n829_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n866_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n868_), .A2(new_n872_), .A3(new_n873_), .ZN(G1343gat));
  INV_X1    g673(.A(new_n861_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n350_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n648_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n279_), .A3(new_n719_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G141gat), .B1(new_n877_), .B2(new_n572_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n280_), .A3(new_n268_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G148gat), .B1(new_n877_), .B2(new_n267_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1345gat));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n878_), .B2(new_n642_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n885_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n877_), .A2(new_n633_), .A3(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1346gat));
  NOR3_X1   g688(.A1(new_n877_), .A2(new_n602_), .A3(new_n677_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n878_), .A2(new_n869_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n602_), .B2(new_n891_), .ZN(G1347gat));
  NOR3_X1   g691(.A1(new_n648_), .A2(new_n349_), .A3(new_n534_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n845_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n719_), .A2(new_n386_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT124), .Z(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n845_), .A2(new_n719_), .A3(new_n893_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(G169gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n899_), .B2(G169gat), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n902_), .A2(new_n903_), .A3(KEYINPUT62), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n899_), .A2(G169gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT123), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n907_), .B2(new_n901_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n898_), .B1(new_n904_), .B2(new_n908_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n895_), .B2(new_n268_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n861_), .A2(new_n387_), .A3(new_n267_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n893_), .B2(new_n911_), .ZN(G1349gat));
  AOI21_X1  g711(.A(G183gat), .B1(new_n862_), .B2(new_n893_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n894_), .A2(new_n633_), .A3(new_n411_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n894_), .B2(new_n677_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n869_), .A2(new_n410_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n894_), .B2(new_n917_), .ZN(G1351gat));
  NOR2_X1   g717(.A1(new_n581_), .A2(new_n531_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n826_), .A2(new_n650_), .A3(new_n828_), .A4(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(G197gat), .A3(new_n719_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n921_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n719_), .ZN(new_n925_));
  INV_X1    g724(.A(G197gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n920_), .B2(new_n572_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT126), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n929_), .B(new_n926_), .C1(new_n920_), .C2(new_n572_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n924_), .A2(new_n925_), .B1(new_n928_), .B2(new_n930_), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n920_), .A2(new_n267_), .ZN(new_n932_));
  XOR2_X1   g731(.A(KEYINPUT127), .B(G204gat), .Z(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1353gat));
  NAND2_X1  g733(.A1(new_n921_), .A2(new_n642_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT63), .B(G211gat), .Z(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n920_), .A2(new_n939_), .A3(new_n677_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n921_), .A2(new_n869_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n939_), .ZN(G1355gat));
endmodule


