//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT10), .B(G99gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G85gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G92gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n220_));
  OAI22_X1  g019(.A1(KEYINPUT9), .A2(new_n216_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n212_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n219_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n225_), .B1(new_n229_), .B2(new_n210_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n223_), .A2(new_n219_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n207_), .A2(new_n209_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n226_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n234_), .B(new_n232_), .C1(new_n235_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT67), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n233_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n244_), .B(new_n225_), .C1(new_n229_), .C2(new_n210_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n226_), .B(new_n239_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n248_), .B2(new_n234_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n245_), .A2(new_n249_), .A3(new_n232_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n243_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT8), .B1(new_n230_), .B2(KEYINPUT68), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n253_), .B2(new_n245_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n224_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G29gat), .B(G36gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G43gat), .B(G50gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT74), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT76), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n262_), .A2(new_n264_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT75), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n266_), .B2(new_n265_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n233_), .A2(new_n242_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n248_), .A2(new_n234_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n244_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n248_), .A2(KEYINPUT68), .A3(new_n234_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n273_), .A2(new_n251_), .A3(KEYINPUT8), .A4(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n254_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n212_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT9), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n213_), .A2(new_n214_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n217_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT64), .ZN(new_n281_));
  INV_X1    g080(.A(new_n220_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n278_), .A2(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n277_), .B1(new_n283_), .B2(new_n222_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n276_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n258_), .B(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n270_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n260_), .A2(new_n267_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n267_), .B1(new_n260_), .B2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n205_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n204_), .B(KEYINPUT36), .Z(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(new_n295_), .A3(KEYINPUT37), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n292_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n293_), .A2(KEYINPUT77), .A3(new_n289_), .A4(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n300_), .B2(KEYINPUT37), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G57gat), .B(G64gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT11), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(KEYINPUT11), .ZN(new_n304_));
  XOR2_X1   g103(.A(G71gat), .B(G78gat), .Z(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n304_), .A2(new_n305_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G231gat), .A2(G233gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n308_), .B(new_n309_), .Z(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G8gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT78), .ZN(new_n312_));
  INV_X1    g111(.A(G15gat), .ZN(new_n313_));
  INV_X1    g112(.A(G22gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G15gat), .A2(G22gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G1gat), .A2(G8gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n315_), .A2(new_n316_), .B1(KEYINPUT14), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n312_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n310_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G127gat), .B(G155gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G183gat), .B(G211gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT17), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n320_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT80), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n325_), .A2(new_n326_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n320_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n301_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n255_), .A2(new_n308_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n276_), .A2(new_n308_), .A3(new_n284_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n336_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(KEYINPUT70), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT71), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n308_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n285_), .A2(new_n345_), .B1(KEYINPUT71), .B2(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(KEYINPUT71), .ZN(new_n347_));
  AOI211_X1 g146(.A(new_n308_), .B(new_n347_), .C1(new_n276_), .C2(new_n284_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n344_), .B(new_n335_), .C1(new_n346_), .C2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n340_), .A2(KEYINPUT70), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G120gat), .B(G148gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT5), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G176gat), .B(G204gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n351_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT13), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT26), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT84), .Z(new_n363_));
  OR2_X1    g162(.A1(new_n361_), .A2(KEYINPUT26), .ZN(new_n364_));
  INV_X1    g163(.A(G183gat), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n365_), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT25), .B1(new_n365_), .B2(KEYINPUT83), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n363_), .A2(new_n364_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n369_), .A2(KEYINPUT24), .A3(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(KEYINPUT85), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(KEYINPUT24), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(G183gat), .A3(G190gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT86), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT23), .B1(new_n365_), .B2(new_n361_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n371_), .A2(KEYINPUT85), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n368_), .A2(new_n374_), .A3(new_n379_), .A4(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(G176gat), .B1(KEYINPUT87), .B2(KEYINPUT22), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G169gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n376_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT30), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT89), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(KEYINPUT89), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  INV_X1    g191(.A(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT88), .B(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  MUX2_X1   g197(.A(new_n390_), .B(new_n391_), .S(new_n398_), .Z(new_n399_));
  XOR2_X1   g198(.A(G127gat), .B(G134gat), .Z(new_n400_));
  XOR2_X1   g199(.A(G113gat), .B(G120gat), .Z(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT31), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n399_), .B(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G155gat), .B(G162gat), .Z(new_n409_));
  INV_X1    g208(.A(KEYINPUT1), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n405_), .A2(KEYINPUT91), .A3(KEYINPUT3), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT3), .B1(new_n405_), .B2(KEYINPUT91), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n407_), .A2(KEYINPUT92), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT2), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n409_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT28), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G22gat), .B(G50gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT96), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n427_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n420_), .A2(new_n421_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G211gat), .B(G218gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G197gat), .B(G204gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT21), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(new_n434_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n432_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(new_n432_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT95), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT93), .Z(new_n442_));
  OR3_X1    g241(.A1(new_n431_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT94), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n439_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n442_), .B1(new_n431_), .B2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n430_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n428_), .A2(new_n448_), .A3(new_n429_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT20), .B1(new_n445_), .B2(new_n388_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT97), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n453_), .A2(new_n454_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G169gat), .ZN(new_n457_));
  INV_X1    g256(.A(G176gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n379_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n370_), .B(new_n459_), .C1(new_n460_), .C2(new_n386_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT99), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(KEYINPUT25), .B(G183gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT98), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n364_), .A2(new_n362_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n385_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n439_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n455_), .A2(new_n456_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G226gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT19), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n463_), .A2(new_n439_), .A3(new_n469_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n476_), .A2(KEYINPUT100), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n445_), .B2(new_n388_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n476_), .B2(KEYINPUT100), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n475_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G8gat), .B(G36gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G64gat), .B(G92gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n482_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n413_), .A2(new_n419_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(new_n402_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT4), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n491_), .A3(new_n402_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G225gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT102), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n490_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n493_), .A2(new_n497_), .B1(new_n498_), .B2(new_n495_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G1gat), .B(G29gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(G85gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT0), .B(G57gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(KEYINPUT103), .A3(KEYINPUT33), .ZN(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT104), .B(KEYINPUT33), .Z(new_n507_));
  OR2_X1    g306(.A1(new_n490_), .A2(KEYINPUT105), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n490_), .A2(KEYINPUT105), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n496_), .A3(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n494_), .A2(new_n495_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n503_), .B1(new_n493_), .B2(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n504_), .A2(new_n507_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT103), .B1(new_n505_), .B2(KEYINPUT33), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n488_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n487_), .A2(KEYINPUT32), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n482_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT106), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n499_), .A2(new_n503_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n505_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n471_), .A2(new_n475_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n479_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n440_), .A2(new_n469_), .A3(new_n461_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n473_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(KEYINPUT32), .A3(new_n487_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(new_n522_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n452_), .B1(new_n516_), .B2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n450_), .A2(new_n521_), .A3(new_n451_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT107), .B(KEYINPUT27), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n488_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n482_), .A2(new_n487_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n487_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n536_), .A3(KEYINPUT27), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n531_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n404_), .B1(new_n530_), .B2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n533_), .A2(new_n537_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n452_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n404_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n522_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT108), .ZN(new_n545_));
  INV_X1    g344(.A(new_n258_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n286_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n319_), .B(new_n546_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(new_n286_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT81), .ZN(new_n551_));
  AND2_X1   g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n549_), .A2(new_n551_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G113gat), .B(G141gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G169gat), .B(G197gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT82), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n553_), .A2(new_n556_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n544_), .A2(new_n545_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n545_), .B1(new_n544_), .B2(new_n560_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n334_), .B(new_n360_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n521_), .B(KEYINPUT109), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n564_), .A2(G1gat), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT38), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n360_), .A2(new_n560_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT110), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n300_), .A2(new_n333_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n544_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(G1gat), .B1(new_n573_), .B2(new_n521_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n569_), .A3(new_n574_), .ZN(G1324gat));
  INV_X1    g374(.A(KEYINPUT111), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n540_), .A2(G8gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n564_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n360_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n544_), .A2(new_n560_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT108), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n582_), .B2(new_n561_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n583_), .A2(KEYINPUT111), .A3(new_n334_), .A4(new_n577_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G8gat), .B1(new_n573_), .B2(new_n540_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT112), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n586_), .A2(new_n587_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n587_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(KEYINPUT39), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n585_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n585_), .A2(KEYINPUT40), .A3(new_n589_), .A4(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1325gat));
  OAI21_X1  g396(.A(G15gat), .B1(new_n573_), .B2(new_n404_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT113), .B(KEYINPUT41), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n542_), .A2(new_n313_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n564_), .B2(new_n601_), .ZN(G1326gat));
  OAI21_X1  g401(.A(G22gat), .B1(new_n573_), .B2(new_n541_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT42), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n452_), .A2(new_n314_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n604_), .B1(new_n564_), .B2(new_n605_), .ZN(G1327gat));
  INV_X1    g405(.A(new_n300_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(new_n332_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n360_), .B(new_n608_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(G29gat), .B1(new_n610_), .B2(new_n522_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n571_), .A2(new_n333_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n544_), .A2(new_n613_), .A3(new_n301_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n544_), .B2(new_n301_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT44), .B(new_n612_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n565_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(G29gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n611_), .B1(new_n620_), .B2(new_n622_), .ZN(G1328gat));
  INV_X1    g422(.A(new_n540_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(new_n624_), .A3(new_n619_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G36gat), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n540_), .A2(G36gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT45), .B1(new_n609_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT45), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n583_), .A2(new_n630_), .A3(new_n608_), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT46), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n626_), .A2(KEYINPUT46), .A3(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1329gat));
  NAND4_X1  g436(.A1(new_n618_), .A2(G43gat), .A3(new_n542_), .A4(new_n619_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n393_), .B1(new_n609_), .B2(new_n404_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g440(.A(G50gat), .B1(new_n610_), .B2(new_n452_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n452_), .A2(G50gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n620_), .B2(new_n643_), .ZN(G1331gat));
  NOR2_X1   g443(.A1(new_n360_), .A2(new_n560_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n544_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(new_n572_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G57gat), .B1(new_n648_), .B2(new_n521_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n646_), .A2(new_n334_), .ZN(new_n650_));
  INV_X1    g449(.A(G57gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n621_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(G1332gat));
  INV_X1    g452(.A(G64gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n647_), .B2(new_n624_), .ZN(new_n655_));
  XOR2_X1   g454(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n650_), .A2(new_n654_), .A3(new_n624_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1333gat));
  INV_X1    g458(.A(G71gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n647_), .B2(new_n542_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT49), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n650_), .A2(new_n660_), .A3(new_n542_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1334gat));
  INV_X1    g463(.A(G78gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n452_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT115), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n650_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT50), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n647_), .A2(new_n452_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(G78gat), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT50), .B(new_n665_), .C1(new_n647_), .C2(new_n452_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT116), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT116), .B(new_n668_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1335gat));
  NAND2_X1  g476(.A1(new_n646_), .A2(new_n608_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G85gat), .B1(new_n679_), .B2(new_n621_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n614_), .A2(new_n615_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n645_), .A2(new_n333_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n521_), .A2(new_n213_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1336gat));
  AOI21_X1  g484(.A(G92gat), .B1(new_n679_), .B2(new_n624_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n540_), .A2(new_n214_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n683_), .B2(new_n687_), .ZN(G1337gat));
  NOR3_X1   g487(.A1(new_n678_), .A2(new_n211_), .A3(new_n404_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n683_), .A2(new_n542_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G99gat), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT51), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(G1338gat));
  NAND3_X1  g492(.A1(new_n679_), .A2(new_n238_), .A3(new_n452_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n682_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n452_), .B(new_n695_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT52), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(G106gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G106gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g500(.A1(new_n543_), .A2(new_n565_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n351_), .A2(new_n355_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT55), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n349_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n347_), .B1(new_n255_), .B2(new_n308_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n285_), .A2(KEYINPUT71), .A3(new_n342_), .A4(new_n345_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n708_), .A2(KEYINPUT55), .A3(new_n335_), .A4(new_n344_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n344_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n336_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT117), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n705_), .A2(new_n709_), .A3(KEYINPUT117), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT56), .B1(new_n716_), .B2(new_n355_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  INV_X1    g517(.A(new_n355_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n718_), .B(new_n719_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n703_), .B(new_n560_), .C1(new_n717_), .C2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n551_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n549_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n556_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n553_), .A2(new_n556_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n356_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n721_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n607_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT118), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n300_), .B1(new_n721_), .B2(new_n726_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT118), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(KEYINPUT57), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n719_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT56), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT58), .A3(new_n703_), .A4(new_n725_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n703_), .B(new_n725_), .C1(new_n717_), .C2(new_n720_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT58), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n741_), .A3(new_n301_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n735_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n332_), .B1(new_n734_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n560_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n334_), .A2(new_n360_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n702_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G113gat), .B1(new_n750_), .B2(new_n560_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT120), .ZN(new_n752_));
  INV_X1    g551(.A(new_n748_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n733_), .B1(new_n731_), .B2(KEYINPUT118), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n729_), .B(new_n300_), .C1(new_n721_), .C2(new_n726_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n735_), .B(new_n742_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n756_), .A2(KEYINPUT121), .A3(new_n333_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT121), .B1(new_n756_), .B2(new_n333_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n702_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(KEYINPUT59), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n759_), .A2(new_n761_), .B1(KEYINPUT59), .B2(new_n749_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n762_), .A2(G113gat), .A3(new_n560_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n752_), .A2(new_n763_), .ZN(G1340gat));
  INV_X1    g563(.A(KEYINPUT123), .ZN(new_n765_));
  INV_X1    g564(.A(G120gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n762_), .B2(new_n580_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT60), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n360_), .A2(KEYINPUT60), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n766_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT122), .B1(new_n750_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT122), .ZN(new_n772_));
  INV_X1    g571(.A(new_n770_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n749_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n765_), .B1(new_n767_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n749_), .A2(KEYINPUT59), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n744_), .A2(KEYINPUT121), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n756_), .A2(new_n333_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT121), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n748_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n761_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n580_), .B(new_n777_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G120gat), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n749_), .A2(new_n773_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT122), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n787_), .A3(KEYINPUT123), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n776_), .A2(new_n788_), .ZN(G1341gat));
  INV_X1    g588(.A(G127gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n762_), .B2(new_n332_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n749_), .A2(G127gat), .A3(new_n333_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1342gat));
  INV_X1    g592(.A(G134gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n750_), .A2(new_n794_), .A3(new_n300_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n762_), .A2(new_n301_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n794_), .ZN(G1343gat));
  NOR2_X1   g596(.A1(new_n744_), .A2(new_n748_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(new_n542_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n624_), .A2(new_n565_), .A3(new_n541_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n745_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT124), .B(G141gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1344gat));
  NOR2_X1   g603(.A1(new_n801_), .A2(new_n360_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT125), .B(G148gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1345gat));
  NOR2_X1   g606(.A1(new_n801_), .A2(new_n333_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT61), .B(G155gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  AND3_X1   g609(.A1(new_n799_), .A2(new_n301_), .A3(new_n800_), .ZN(new_n811_));
  INV_X1    g610(.A(G162gat), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n300_), .A2(new_n812_), .ZN(new_n813_));
  OAI22_X1  g612(.A1(new_n811_), .A2(new_n812_), .B1(new_n801_), .B2(new_n813_), .ZN(G1347gat));
  NOR3_X1   g613(.A1(new_n540_), .A2(new_n621_), .A3(new_n404_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n452_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n759_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n560_), .A3(new_n457_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n759_), .A2(new_n560_), .A3(new_n817_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT62), .B1(new_n820_), .B2(G169gat), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1348gat));
  AOI21_X1  g623(.A(G176gat), .B1(new_n818_), .B2(new_n580_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n798_), .A2(new_n452_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n816_), .A2(new_n458_), .A3(new_n360_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(G1349gat));
  NOR4_X1   g627(.A1(new_n798_), .A2(new_n333_), .A3(new_n452_), .A4(new_n816_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n829_), .A2(KEYINPUT126), .ZN(new_n830_));
  AOI21_X1  g629(.A(G183gat), .B1(new_n829_), .B2(KEYINPUT126), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n333_), .A2(new_n465_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n830_), .A2(new_n831_), .B1(new_n818_), .B2(new_n832_), .ZN(G1350gat));
  NAND3_X1  g632(.A1(new_n818_), .A2(new_n300_), .A3(new_n466_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n818_), .A2(new_n301_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n361_), .ZN(G1351gat));
  NOR3_X1   g635(.A1(new_n540_), .A2(new_n541_), .A3(new_n522_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n799_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n560_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n360_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT127), .B(G204gat), .Z(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n842_), .B2(new_n845_), .ZN(G1353gat));
  AOI211_X1 g645(.A(KEYINPUT63), .B(G211gat), .C1(new_n839_), .C2(new_n332_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT63), .B(G211gat), .Z(new_n848_));
  AND3_X1   g647(.A1(new_n839_), .A2(new_n332_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1354gat));
  INV_X1    g649(.A(G218gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n839_), .A2(new_n851_), .A3(new_n300_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n839_), .A2(new_n301_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1355gat));
endmodule


