//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT71), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(KEYINPUT71), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT71), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G1gat), .B(G8gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n210_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n219_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n210_), .B(new_n219_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n220_), .A2(new_n225_), .B1(new_n226_), .B2(new_n222_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G113gat), .B(G141gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(G169gat), .B(G197gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n227_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT23), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT26), .B(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(G183gat), .ZN(new_n243_));
  INV_X1    g042(.A(G183gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT25), .B1(new_n244_), .B2(KEYINPUT77), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n235_), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n237_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n239_), .B1(new_n250_), .B2(KEYINPUT78), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n252_), .A3(new_n249_), .ZN(new_n253_));
  OR2_X1    g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n234_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT79), .B(G176gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT22), .B(G169gat), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n256_), .A2(new_n257_), .B1(G169gat), .B2(G176gat), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n251_), .A2(new_n253_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(G15gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n259_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT31), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G43gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT81), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n271_));
  INV_X1    g070(.A(G127gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(G134gat), .ZN(new_n273_));
  INV_X1    g072(.A(G134gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(G127gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G113gat), .B(G120gat), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n270_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n268_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n264_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n234_), .A2(new_n238_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT25), .B(G183gat), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n240_), .A2(new_n286_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n285_), .A2(new_n287_), .B1(new_n258_), .B2(new_n255_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G197gat), .A2(G204gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT88), .B(G204gat), .ZN(new_n291_));
  INV_X1    g090(.A(G197gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  INV_X1    g093(.A(G218gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G211gat), .ZN(new_n296_));
  INV_X1    g095(.A(G211gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G218gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n293_), .A2(new_n294_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G204gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT88), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G204gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n292_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n294_), .B1(new_n307_), .B2(new_n289_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n306_), .A3(new_n292_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n294_), .B1(G197gat), .B2(G204gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n299_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n309_), .B1(new_n308_), .B2(new_n312_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n288_), .B(new_n302_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n312_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT89), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n301_), .B1(new_n318_), .B2(new_n313_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n316_), .B(KEYINPUT20), .C1(new_n319_), .C2(new_n259_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT19), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT90), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT20), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n319_), .B2(new_n288_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT90), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n251_), .A2(new_n253_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n258_), .A2(new_n255_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n302_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n322_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n325_), .A2(new_n326_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT20), .B1(new_n319_), .B2(new_n288_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n329_), .A2(new_n330_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n322_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n323_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n323_), .A2(new_n336_), .A3(new_n341_), .A4(new_n333_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(KEYINPUT27), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n325_), .A2(new_n322_), .A3(new_n331_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n341_), .B(KEYINPUT96), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT27), .A3(new_n344_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(KEYINPUT1), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(KEYINPUT82), .B(new_n355_), .C1(new_n356_), .C2(KEYINPUT1), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n355_), .A2(new_n361_), .A3(KEYINPUT1), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n355_), .B2(KEYINPUT1), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n359_), .A2(new_n360_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G141gat), .ZN(new_n365_));
  INV_X1    g164(.A(G148gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT3), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT85), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT2), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n371_), .A2(new_n377_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT2), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n368_), .A2(new_n374_), .A3(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n373_), .A2(new_n376_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  XOR2_X1   g181(.A(G155gat), .B(G162gat), .Z(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n370_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n281_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT91), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n280_), .B(new_n370_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n281_), .A3(KEYINPUT91), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT4), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n386_), .A2(new_n394_), .A3(new_n281_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n401_));
  AOI211_X1 g200(.A(KEYINPUT92), .B(new_n397_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n399_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n399_), .B(new_n407_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n386_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT28), .Z(new_n416_));
  OAI21_X1  g215(.A(new_n330_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n417_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G228gat), .ZN(new_n421_));
  INV_X1    g220(.A(G233gat), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT87), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(KEYINPUT87), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G78gat), .ZN(new_n426_));
  INV_X1    g225(.A(G106gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n420_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n418_), .A2(new_n419_), .A3(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n354_), .A2(new_n412_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n349_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n337_), .B2(new_n437_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n410_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n392_), .A2(new_n396_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT92), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n392_), .A2(new_n400_), .A3(new_n396_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(KEYINPUT33), .A3(new_n399_), .A4(new_n407_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n394_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n395_), .A2(new_n396_), .ZN(new_n449_));
  OR3_X1    g248(.A1(new_n448_), .A2(KEYINPUT93), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT93), .B1(new_n448_), .B2(new_n449_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n407_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n442_), .A2(new_n447_), .A3(new_n345_), .A4(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n440_), .B1(new_n454_), .B2(KEYINPUT94), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n343_), .A2(new_n344_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n451_), .A2(new_n452_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n447_), .A4(new_n442_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n434_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n435_), .B1(new_n461_), .B2(KEYINPUT95), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT95), .ZN(new_n463_));
  AOI211_X1 g262(.A(new_n463_), .B(new_n434_), .C1(new_n455_), .C2(new_n460_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n284_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n353_), .A2(new_n434_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n412_), .A3(new_n283_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT97), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT97), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n466_), .A2(new_n469_), .A3(new_n412_), .A4(new_n283_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n232_), .B1(new_n465_), .B2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n427_), .A3(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT9), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n477_), .A2(KEYINPUT9), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n475_), .A2(new_n478_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT65), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n489_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n481_), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n486_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n480_), .A2(new_n482_), .B1(new_n493_), .B2(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n488_), .A2(new_n490_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT66), .ZN(new_n501_));
  AND2_X1   g300(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n502_));
  NOR2_X1   g301(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G85gat), .B(G92gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n499_), .A2(new_n500_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n505_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT8), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n508_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n509_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n485_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G71gat), .B(G78gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G64gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G57gat), .ZN(new_n519_));
  INV_X1    g318(.A(G57gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G64gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n521_), .A3(KEYINPUT11), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n516_), .B1(KEYINPUT11), .B2(new_n524_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT12), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n527_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT66), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT66), .B1(new_n499_), .B2(new_n500_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n506_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n510_), .B2(new_n505_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n485_), .B(new_n530_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT12), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n506_), .B1(new_n510_), .B2(new_n486_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n501_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n485_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n527_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n515_), .A2(new_n529_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G230gat), .A2(G233gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT64), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n540_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(new_n530_), .ZN(new_n548_));
  AOI211_X1 g347(.A(new_n540_), .B(new_n527_), .C1(new_n508_), .C2(new_n512_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G120gat), .B(G148gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n545_), .A2(new_n550_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(KEYINPUT70), .A3(new_n559_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT13), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(KEYINPUT13), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n212_), .A2(new_n515_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT34), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n223_), .B2(new_n547_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT36), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n578_), .B(KEYINPUT36), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n581_), .B(KEYINPUT73), .Z(new_n587_));
  NOR2_X1   g386(.A1(new_n575_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT37), .B1(new_n580_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n527_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT75), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n219_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n594_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n590_), .A2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n472_), .A2(new_n567_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n214_), .A3(new_n411_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT38), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n567_), .A2(new_n231_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n465_), .A2(new_n471_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n584_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT98), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT98), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n610_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n411_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n618_), .A2(KEYINPUT99), .A3(G1gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT99), .B1(new_n618_), .B2(G1gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n608_), .B1(new_n619_), .B2(new_n620_), .ZN(G1324gat));
  NAND3_X1  g420(.A1(new_n606_), .A2(new_n215_), .A3(new_n353_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n353_), .B(new_n610_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n623_), .A2(new_n624_), .A3(G8gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n623_), .B2(G8gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(KEYINPUT40), .B(new_n622_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n616_), .B2(new_n284_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n634_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n606_), .A2(new_n261_), .A3(new_n283_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n606_), .A2(new_n639_), .A3(new_n434_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n617_), .A2(new_n434_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(G22gat), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT42), .B(new_n639_), .C1(new_n617_), .C2(new_n434_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(G1327gat));
  INV_X1    g444(.A(new_n604_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n612_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n567_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n472_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n411_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n586_), .A2(new_n589_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(KEYINPUT43), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n432_), .A2(new_n433_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n353_), .A2(new_n654_), .A3(new_n411_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n454_), .A2(KEYINPUT94), .ZN(new_n656_));
  INV_X1    g455(.A(new_n440_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n460_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n654_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n655_), .B1(new_n659_), .B2(new_n463_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n461_), .A2(KEYINPUT95), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n283_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n468_), .A2(new_n470_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n653_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n652_), .B(KEYINPUT102), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n465_), .B2(new_n471_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n609_), .A2(new_n646_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(KEYINPUT44), .A3(new_n670_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n411_), .A2(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n651_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  NAND3_X1  g476(.A1(new_n673_), .A2(new_n353_), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G36gat), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n649_), .A2(G36gat), .A3(new_n354_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT45), .Z(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(KEYINPUT103), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT103), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(new_n681_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1329gat));
  NAND4_X1  g486(.A1(new_n673_), .A2(G43gat), .A3(new_n283_), .A4(new_n674_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n649_), .A2(new_n284_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(G43gat), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g490(.A(G50gat), .B1(new_n650_), .B2(new_n434_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n434_), .A2(G50gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n675_), .B2(new_n693_), .ZN(G1331gat));
  INV_X1    g493(.A(new_n567_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n232_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n465_), .B2(new_n471_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(new_n605_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n520_), .A3(new_n411_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n614_), .A2(new_n615_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n700_), .A2(new_n604_), .A3(new_n696_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n411_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n702_), .B2(new_n520_), .ZN(G1332gat));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n518_), .A3(new_n353_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n353_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(G64gat), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT48), .B(new_n518_), .C1(new_n701_), .C2(new_n353_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1333gat));
  INV_X1    g508(.A(G71gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n698_), .A2(new_n710_), .A3(new_n283_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT49), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n701_), .A2(new_n283_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(G71gat), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT49), .B(new_n710_), .C1(new_n701_), .C2(new_n283_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(G1334gat));
  INV_X1    g515(.A(G78gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n698_), .A2(new_n717_), .A3(new_n434_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n701_), .A2(new_n434_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G78gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT50), .B(new_n717_), .C1(new_n701_), .C2(new_n434_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1335gat));
  AND2_X1   g522(.A1(new_n697_), .A2(new_n647_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n411_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n696_), .A2(new_n646_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n669_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n411_), .A2(G85gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT104), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n728_), .B2(new_n730_), .ZN(G1336gat));
  OAI21_X1  g530(.A(G92gat), .B1(new_n727_), .B2(new_n354_), .ZN(new_n732_));
  INV_X1    g531(.A(G92gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n733_), .A3(new_n353_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1337gat));
  OAI21_X1  g534(.A(G99gat), .B1(new_n727_), .B2(new_n284_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n724_), .A2(new_n473_), .A3(new_n474_), .A4(new_n283_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g538(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n669_), .A2(new_n434_), .A3(new_n726_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT106), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n669_), .A2(new_n744_), .A3(new_n434_), .A4(new_n726_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n743_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n697_), .A2(new_n427_), .A3(new_n434_), .A4(new_n647_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT105), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n745_), .A2(G106gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT52), .B1(new_n750_), .B2(new_n743_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n741_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  INV_X1    g552(.A(new_n743_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n745_), .A2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n756_), .A2(new_n746_), .A3(new_n748_), .A4(new_n740_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n752_), .A2(new_n757_), .ZN(G1339gat));
  NOR2_X1   g557(.A1(new_n412_), .A2(new_n284_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n466_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n231_), .A2(new_n559_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT110), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT68), .B1(new_n533_), .B2(new_n535_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n508_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n540_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT12), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n547_), .B2(new_n530_), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n768_), .A2(new_n528_), .B1(new_n770_), .B2(new_n548_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n546_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n515_), .A2(new_n529_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n541_), .B1(new_n549_), .B2(new_n769_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n544_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT55), .B1(new_n542_), .B2(new_n544_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT111), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n771_), .B2(new_n546_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n772_), .A4(new_n775_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n558_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n765_), .B1(new_n783_), .B2(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n783_), .A2(new_n765_), .A3(KEYINPUT56), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n764_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n220_), .B(new_n222_), .C1(new_n210_), .C2(new_n219_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n230_), .B1(new_n226_), .B2(new_n221_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n789_), .A2(new_n790_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n562_), .A2(new_n563_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n584_), .B1(new_n788_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n762_), .B1(new_n794_), .B2(KEYINPUT57), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n778_), .A2(new_n782_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT112), .B(new_n796_), .C1(new_n797_), .C2(new_n558_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n785_), .A3(new_n784_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n792_), .B1(new_n799_), .B2(new_n764_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  NOR4_X1   g600(.A1(new_n800_), .A2(KEYINPUT115), .A3(new_n801_), .A4(new_n584_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n795_), .A2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n791_), .A2(new_n559_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n783_), .A2(KEYINPUT56), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n796_), .B(new_n558_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n804_), .B(KEYINPUT113), .C1(new_n805_), .C2(new_n806_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n804_), .B(KEYINPUT58), .C1(new_n805_), .C2(new_n806_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n652_), .B1(new_n813_), .B2(KEYINPUT114), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(KEYINPUT114), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n801_), .B1(new_n800_), .B2(new_n584_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n761_), .B1(new_n803_), .B2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n816_), .A2(new_n817_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(KEYINPUT116), .C1(new_n795_), .C2(new_n802_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n604_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n605_), .A2(new_n567_), .A3(new_n232_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT109), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OR3_X1    g625(.A1(new_n823_), .A2(new_n824_), .A3(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n824_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n826_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n760_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n231_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(KEYINPUT117), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(KEYINPUT117), .ZN(new_n834_));
  INV_X1    g633(.A(new_n830_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n817_), .B(new_n816_), .C1(new_n795_), .C2(new_n802_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n646_), .B1(new_n836_), .B2(new_n761_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n821_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT59), .B1(new_n838_), .B2(new_n760_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n760_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n836_), .A2(new_n604_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n840_), .B(new_n841_), .C1(new_n842_), .C2(new_n835_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n839_), .A2(new_n843_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT119), .B(G113gat), .Z(new_n845_));
  NOR2_X1   g644(.A1(new_n232_), .A2(new_n845_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n833_), .A2(new_n834_), .B1(new_n844_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n695_), .B(new_n843_), .C1(new_n831_), .C2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT120), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n839_), .A2(new_n851_), .A3(new_n695_), .A4(new_n843_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(G120gat), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n567_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n831_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n831_), .A2(new_n272_), .A3(new_n646_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n839_), .A2(new_n646_), .A3(new_n843_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n860_), .B2(new_n272_), .ZN(G1342gat));
  NAND3_X1  g660(.A1(new_n831_), .A2(new_n274_), .A3(new_n584_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n839_), .A2(new_n590_), .A3(new_n843_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n864_), .B2(new_n274_), .ZN(G1343gat));
  NOR2_X1   g664(.A1(new_n654_), .A2(new_n283_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n867_), .A2(new_n353_), .A3(new_n412_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n231_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n695_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT121), .B(G148gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1345gat));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n870_), .A2(new_n876_), .A3(new_n646_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n870_), .B2(new_n646_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n878_), .A2(new_n879_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n870_), .A2(new_n646_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT122), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n880_), .B1(new_n884_), .B2(new_n877_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n885_), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n870_), .B2(new_n584_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n665_), .A2(G162gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n870_), .B2(new_n888_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n842_), .A2(new_n835_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n353_), .A2(new_n412_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n284_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n231_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT123), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n654_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n890_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT62), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n842_), .A2(new_n835_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n892_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n434_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n231_), .A2(new_n257_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT124), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n897_), .B1(new_n901_), .B2(new_n903_), .ZN(G1348gat));
  INV_X1    g703(.A(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n695_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n838_), .A2(new_n434_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n567_), .A2(new_n899_), .A3(new_n237_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(new_n256_), .B1(new_n907_), .B2(new_n908_), .ZN(G1349gat));
  NOR2_X1   g708(.A1(new_n604_), .A2(new_n286_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n898_), .A2(new_n900_), .A3(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT125), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n899_), .A2(new_n604_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G183gat), .B1(new_n907_), .B2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n901_), .B2(new_n652_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n584_), .A2(new_n240_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n901_), .B2(new_n917_), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n822_), .A2(new_n830_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n867_), .A2(new_n891_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n232_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n292_), .ZN(G1352gat));
  INV_X1    g722(.A(new_n921_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(KEYINPUT126), .A3(new_n695_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n921_), .B2(new_n567_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(G204gat), .A3(new_n927_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n919_), .A2(new_n291_), .A3(new_n695_), .A4(new_n920_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n928_), .A2(new_n931_), .ZN(G1353gat));
  AOI211_X1 g731(.A(KEYINPUT63), .B(G211gat), .C1(new_n924_), .C2(new_n646_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT63), .B(G211gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n921_), .A2(new_n604_), .A3(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1354gat));
  OAI21_X1  g735(.A(G218gat), .B1(new_n921_), .B2(new_n652_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n584_), .A2(new_n295_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n921_), .B2(new_n938_), .ZN(G1355gat));
endmodule


