//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n982_, new_n983_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1008_, new_n1009_, new_n1010_, new_n1012_, new_n1013_, new_n1015_,
    new_n1016_, new_n1017_, new_n1019_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1033_, new_n1034_, new_n1035_;
  INV_X1    g000(.A(KEYINPUT106), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT93), .ZN(new_n203_));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT93), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(KEYINPUT92), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n212_), .B(new_n213_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n206_), .B(new_n209_), .C1(new_n216_), .C2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n208_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n210_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n217_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n207_), .A2(new_n222_), .A3(new_n208_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G127gat), .B(G134gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n209_), .A2(new_n206_), .ZN(new_n233_));
  INV_X1    g032(.A(G141gat), .ZN(new_n234_));
  INV_X1    g033(.A(G148gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n218_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT3), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n237_), .A2(new_n219_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n233_), .A2(new_n238_), .B1(new_n226_), .B2(new_n225_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n229_), .B(new_n230_), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n232_), .A2(new_n241_), .A3(KEYINPUT4), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT4), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n244_), .B(KEYINPUT102), .Z(new_n251_));
  NAND3_X1  g050(.A1(new_n232_), .A2(new_n241_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT33), .B1(new_n245_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n242_), .A2(new_n243_), .A3(new_n251_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n232_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n249_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G8gat), .B(G36gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT18), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT101), .ZN(new_n264_));
  INV_X1    g063(.A(G218gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G211gat), .ZN(new_n266_));
  INV_X1    g065(.A(G211gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G218gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT21), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G197gat), .B(G204gat), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G197gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G204gat), .ZN(new_n275_));
  INV_X1    g074(.A(G204gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G197gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n277_), .A3(KEYINPUT95), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n276_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT96), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .A4(KEYINPUT21), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n269_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n275_), .A2(new_n277_), .A3(KEYINPUT95), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT21), .B1(new_n275_), .B2(KEYINPUT95), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT96), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n273_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT86), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT86), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n293_), .B(new_n288_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n294_));
  AND2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n292_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G183gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT25), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G183gat), .ZN(new_n302_));
  INV_X1    g101(.A(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT26), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G190gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n300_), .A2(new_n302_), .A3(new_n304_), .A4(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT24), .A3(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n307_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n317_));
  NAND2_X1  g116(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n295_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n288_), .A2(KEYINPUT23), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n288_), .A2(KEYINPUT88), .A3(KEYINPUT23), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n299_), .A2(new_n303_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n309_), .A2(KEYINPUT87), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT87), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n308_), .A2(KEYINPUT22), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G169gat), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n327_), .A2(new_n329_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n311_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n298_), .A2(new_n316_), .B1(new_n326_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n264_), .B1(new_n287_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n286_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n273_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n334_), .B1(new_n325_), .B2(new_n324_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n307_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n291_), .A2(KEYINPUT86), .B1(new_n296_), .B2(new_n295_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n294_), .B2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n340_), .B(KEYINPUT101), .C1(new_n341_), .C2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n337_), .A2(new_n345_), .A3(KEYINPUT20), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n334_), .B1(new_n298_), .B2(new_n325_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT100), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n319_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n342_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n300_), .A2(new_n302_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G190gat), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n352_), .A2(new_n353_), .B1(new_n314_), .B2(new_n313_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n354_), .A2(new_n324_), .A3(KEYINPUT100), .A4(new_n312_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n287_), .A2(new_n348_), .A3(new_n351_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT19), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n346_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT20), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n287_), .B2(new_n336_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n343_), .A2(new_n294_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n351_), .B(new_n355_), .C1(new_n364_), .C2(new_n334_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n340_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n359_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n263_), .B1(new_n361_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n326_), .A2(new_n335_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n298_), .A2(new_n316_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n369_), .A2(new_n370_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n362_), .B1(new_n371_), .B2(KEYINPUT101), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(new_n359_), .A3(new_n356_), .A4(new_n337_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n363_), .A2(new_n366_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n358_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n375_), .A3(new_n262_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n255_), .A2(KEYINPUT33), .A3(new_n256_), .A4(new_n249_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n258_), .A2(new_n368_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n350_), .A2(new_n342_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT104), .B1(new_n347_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n316_), .A2(new_n324_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT104), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n381_), .B(new_n382_), .C1(new_n364_), .C2(new_n334_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n380_), .A2(new_n287_), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n358_), .B1(new_n346_), .B2(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n363_), .A2(new_n366_), .A3(new_n359_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n262_), .A2(KEYINPUT32), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n373_), .A2(new_n375_), .A3(KEYINPUT103), .A4(new_n389_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n373_), .A2(new_n375_), .A3(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT103), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n255_), .A2(new_n256_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n250_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT105), .A3(new_n257_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT105), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n400_), .A3(new_n250_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n378_), .B1(new_n396_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n216_), .A2(new_n220_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n209_), .A2(new_n206_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n227_), .B(new_n404_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT28), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT28), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n221_), .A2(new_n409_), .A3(new_n404_), .A4(new_n227_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G22gat), .B(G50gat), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n411_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n409_), .B1(new_n239_), .B2(new_n404_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n410_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT99), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n415_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n423_));
  NAND2_X1  g222(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(G228gat), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n239_), .B2(new_n404_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n423_), .B1(new_n428_), .B2(new_n287_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n404_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n431_), .A2(new_n340_), .A3(KEYINPUT97), .A4(new_n427_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n427_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n340_), .B1(new_n430_), .B2(KEYINPUT98), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n430_), .A2(KEYINPUT98), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G78gat), .B(G106gat), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n433_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n422_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n437_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n438_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n433_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n415_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n399_), .A2(new_n401_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(new_n447_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n376_), .A2(KEYINPUT27), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n262_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT27), .B1(new_n368_), .B2(new_n376_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n403_), .A2(new_n447_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456_));
  INV_X1    g255(.A(G15gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n344_), .B2(new_n341_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n370_), .A2(new_n369_), .A3(new_n459_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n461_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n458_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT90), .B(G43gat), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n344_), .A2(new_n341_), .A3(new_n460_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n459_), .B1(new_n370_), .B2(new_n369_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n462_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n458_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(new_n464_), .A3(new_n463_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n467_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT91), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n468_), .B1(new_n467_), .B2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT31), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n467_), .A2(new_n474_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n468_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT31), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n481_), .A2(KEYINPUT91), .A3(new_n482_), .A4(new_n475_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n478_), .A2(new_n231_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n231_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n202_), .B1(new_n455_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n478_), .A2(new_n483_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n240_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(new_n231_), .A3(new_n483_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n447_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n388_), .A2(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n448_), .A2(new_n493_), .A3(new_n392_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n494_), .B2(new_n378_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n373_), .A2(new_n375_), .A3(new_n262_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n262_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n380_), .A2(new_n287_), .A3(new_n383_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n372_), .A2(new_n337_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n386_), .B1(new_n358_), .B2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(KEYINPUT27), .B(new_n376_), .C1(new_n502_), .C2(new_n262_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n504_), .A2(new_n448_), .A3(new_n447_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n491_), .B(KEYINPUT106), .C1(new_n495_), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n487_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT107), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n447_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n486_), .A2(new_n508_), .A3(new_n402_), .A4(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n489_), .A2(new_n402_), .A3(new_n490_), .A4(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT107), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G169gat), .B(G197gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G8gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT78), .B(G1gat), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n522_), .B2(G8gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(G15gat), .B(G22gat), .Z(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT79), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n523_), .A2(KEYINPUT79), .A3(new_n524_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n520_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(G8gat), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n524_), .B1(new_n529_), .B2(KEYINPUT14), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT79), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n525_), .A3(new_n519_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535_));
  XOR2_X1   g334(.A(G29gat), .B(G36gat), .Z(new_n536_));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G29gat), .B(G36gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT72), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G43gat), .B(G50gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n538_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n536_), .A2(new_n537_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(KEYINPUT72), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n535_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n542_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n545_), .A3(new_n541_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(KEYINPUT15), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n534_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n549_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n528_), .A2(new_n554_), .A3(new_n533_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n526_), .A2(new_n527_), .A3(new_n520_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n519_), .B1(new_n532_), .B2(new_n525_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n553_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n554_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n553_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n555_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT83), .A3(new_n559_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n558_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n518_), .B1(new_n570_), .B2(KEYINPUT84), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT83), .B1(new_n568_), .B2(new_n559_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n565_), .B(new_n556_), .C1(new_n567_), .C2(new_n555_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n557_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT84), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n517_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n514_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT64), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G71gat), .B(G78gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(G57gat), .B(G64gat), .Z(new_n585_));
  INV_X1    g384(.A(KEYINPUT11), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT66), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n590_), .A2(KEYINPUT66), .A3(new_n584_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n583_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n588_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT66), .B1(new_n590_), .B2(new_n584_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT11), .A4(new_n582_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT10), .B(G99gat), .Z(new_n597_));
  INV_X1    g396(.A(G106gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G85gat), .B(G92gat), .Z(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT9), .ZN(new_n601_));
  INV_X1    g400(.A(G85gat), .ZN(new_n602_));
  INV_X1    g401(.A(G92gat), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n602_), .A2(new_n603_), .A3(KEYINPUT9), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT6), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n599_), .A2(new_n601_), .A3(new_n604_), .A4(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n608_));
  OR3_X1    g407(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n606_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT65), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT8), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G85gat), .B(G92gat), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n611_), .B2(KEYINPUT8), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n610_), .B2(new_n614_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n607_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n581_), .B1(new_n596_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n596_), .A2(new_n617_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT12), .B1(new_n620_), .B2(KEYINPUT68), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT68), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n623_));
  AOI211_X1 g422(.A(new_n622_), .B(new_n623_), .C1(new_n596_), .C2(new_n617_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n619_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT67), .B1(new_n596_), .B2(new_n617_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n607_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n610_), .A2(new_n614_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n612_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT67), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n595_), .A4(new_n592_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n634_), .A3(new_n620_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n580_), .ZN(new_n636_));
  XOR2_X1   g435(.A(G120gat), .B(G148gat), .Z(new_n637_));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n639_), .B(new_n640_), .Z(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n625_), .A2(new_n636_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT70), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT70), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n625_), .A2(new_n636_), .A3(new_n645_), .A4(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n630_), .A2(new_n631_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n648_), .A2(new_n607_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n623_), .B1(new_n649_), .B2(new_n622_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n620_), .A2(KEYINPUT68), .A3(KEYINPUT12), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n652_), .A2(new_n619_), .B1(new_n580_), .B2(new_n635_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(new_n642_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n647_), .A2(KEYINPUT13), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT13), .B1(new_n647_), .B2(new_n654_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(G127gat), .B(G155gat), .Z(new_n659_));
  XNOR2_X1  g458(.A(G183gat), .B(G211gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT17), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n664_), .A2(new_n665_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n668_), .B2(KEYINPUT81), .ZN(new_n669_));
  NAND2_X1  g468(.A1(G231gat), .A2(G233gat), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n596_), .B(new_n670_), .Z(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(new_n534_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n665_), .A2(KEYINPUT81), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT82), .B1(new_n663_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n669_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(KEYINPUT82), .B2(new_n667_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n551_), .A2(new_n617_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n632_), .A2(new_n554_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n683_));
  NAND2_X1  g482(.A1(G232gat), .A2(G233gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(KEYINPUT35), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT73), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n551_), .B2(new_n617_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(KEYINPUT35), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n682_), .A2(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n680_), .A2(new_n681_), .A3(new_n687_), .A4(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT76), .ZN(new_n694_));
  XOR2_X1   g493(.A(G190gat), .B(G218gat), .Z(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT74), .ZN(new_n696_));
  XOR2_X1   g495(.A(G134gat), .B(G162gat), .Z(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT36), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT75), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n693_), .A2(new_n694_), .A3(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n698_), .B(KEYINPUT36), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n690_), .A2(new_n703_), .A3(new_n692_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n694_), .B1(new_n693_), .B2(new_n701_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT37), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n704_), .A2(KEYINPUT77), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT37), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n693_), .A2(new_n701_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n704_), .A2(KEYINPUT77), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .A4(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n707_), .A2(new_n712_), .ZN(new_n713_));
  NOR4_X1   g512(.A1(new_n578_), .A2(new_n658_), .A3(new_n679_), .A4(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n402_), .A2(new_n522_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT38), .ZN(new_n717_));
  INV_X1    g516(.A(new_n577_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n658_), .A2(new_n718_), .A3(new_n679_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT108), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n708_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n514_), .A2(KEYINPUT109), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT109), .B1(new_n514_), .B2(new_n721_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G1gat), .B1(new_n724_), .B2(new_n402_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n717_), .A2(new_n725_), .ZN(G1324gat));
  INV_X1    g525(.A(G8gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n714_), .A2(new_n727_), .A3(new_n504_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n720_), .B(new_n504_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT39), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G8gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G8gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT40), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT40), .B(new_n728_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1325gat));
  INV_X1    g536(.A(new_n724_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n457_), .B1(new_n738_), .B2(new_n486_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT41), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n740_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n714_), .A2(new_n457_), .A3(new_n486_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT110), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n741_), .A2(new_n742_), .A3(new_n744_), .ZN(G1326gat));
  INV_X1    g544(.A(G22gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n714_), .A2(new_n746_), .A3(new_n492_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n738_), .A2(new_n492_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G22gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT42), .B(new_n746_), .C1(new_n738_), .C2(new_n492_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1327gat));
  NOR3_X1   g551(.A1(new_n658_), .A2(new_n718_), .A3(new_n678_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n514_), .B2(new_n713_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n707_), .A2(new_n712_), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT43), .B(new_n756_), .C1(new_n507_), .C2(new_n513_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n487_), .A2(new_n506_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n761_), .B2(new_n756_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n514_), .A2(new_n754_), .A3(new_n713_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(KEYINPUT44), .A3(new_n753_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n448_), .A2(G29gat), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n760_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n678_), .A2(new_n721_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n657_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n578_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G29gat), .B1(new_n770_), .B2(new_n448_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n767_), .A2(KEYINPUT111), .A3(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT111), .B1(new_n767_), .B2(new_n771_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1328gat));
  XNOR2_X1  g573(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n760_), .A2(new_n504_), .A3(new_n765_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G36gat), .ZN(new_n777_));
  INV_X1    g576(.A(new_n769_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n454_), .A2(G36gat), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n514_), .A2(new_n577_), .A3(new_n778_), .A4(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT45), .Z(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n775_), .B1(new_n777_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n775_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n781_), .B(new_n784_), .C1(new_n776_), .C2(G36gat), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1329gat));
  AND4_X1   g585(.A1(G43gat), .A2(new_n760_), .A3(new_n486_), .A4(new_n765_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G43gat), .B1(new_n770_), .B2(new_n486_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT47), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n764_), .A2(KEYINPUT44), .A3(new_n753_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT44), .B1(new_n764_), .B2(new_n753_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(G43gat), .A3(new_n486_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n788_), .B(KEYINPUT113), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n791_), .A2(new_n798_), .ZN(G1330gat));
  AOI21_X1  g598(.A(G50gat), .B1(new_n770_), .B2(new_n492_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n492_), .A2(G50gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n794_), .B2(new_n801_), .ZN(G1331gat));
  NOR2_X1   g601(.A1(new_n657_), .A2(new_n577_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n678_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT114), .B(new_n805_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(G57gat), .A3(new_n448_), .A4(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(KEYINPUT115), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(KEYINPUT115), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n761_), .A2(new_n657_), .A3(new_n577_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n713_), .A2(new_n679_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G57gat), .B1(new_n816_), .B2(new_n448_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n811_), .A2(new_n812_), .A3(new_n817_), .ZN(G1332gat));
  OR3_X1    g617(.A1(new_n815_), .A2(G64gat), .A3(new_n454_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n808_), .A2(new_n504_), .A3(new_n809_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT48), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(G64gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(G64gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(G1333gat));
  OR3_X1    g623(.A1(new_n815_), .A2(G71gat), .A3(new_n491_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n808_), .A2(new_n486_), .A3(new_n809_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n826_), .A2(new_n827_), .A3(G71gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(G71gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(G1334gat));
  OR3_X1    g629(.A1(new_n815_), .A2(G78gat), .A3(new_n447_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n808_), .A2(new_n492_), .A3(new_n809_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G78gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G78gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(G1335gat));
  NAND2_X1  g635(.A1(new_n764_), .A2(KEYINPUT116), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n803_), .A2(new_n679_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n762_), .A2(new_n763_), .A3(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n837_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G85gat), .B1(new_n842_), .B2(new_n402_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n813_), .A2(new_n768_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n602_), .A3(new_n448_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1336gat));
  OAI21_X1  g645(.A(G92gat), .B1(new_n842_), .B2(new_n454_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n603_), .A3(new_n504_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1337gat));
  NAND4_X1  g648(.A1(new_n837_), .A2(new_n486_), .A3(new_n839_), .A4(new_n841_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G99gat), .ZN(new_n851_));
  OR2_X1    g650(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n486_), .A2(new_n597_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n844_), .A2(new_n853_), .B1(KEYINPUT117), .B2(KEYINPUT51), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n851_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n852_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1338gat));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n755_), .A2(new_n757_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n839_), .A2(new_n492_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n858_), .B(G106gat), .C1(new_n859_), .C2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n862_), .B2(new_n598_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n863_), .A3(KEYINPUT52), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT118), .B(new_n865_), .C1(new_n862_), .C2(new_n598_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n844_), .A2(new_n598_), .A3(new_n492_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT53), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n864_), .A2(new_n870_), .A3(new_n866_), .A4(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1339gat));
  NAND3_X1  g671(.A1(new_n814_), .A2(new_n657_), .A3(new_n718_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT54), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n814_), .A2(new_n875_), .A3(new_n657_), .A4(new_n718_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n645_), .B1(new_n653_), .B2(new_n642_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n646_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n571_), .B(new_n576_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n626_), .A2(new_n634_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n618_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n882_), .A2(new_n581_), .B1(new_n883_), .B2(KEYINPUT55), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n625_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n641_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n621_), .A2(new_n624_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n580_), .B1(new_n890_), .B2(new_n881_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n625_), .A2(new_n885_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n883_), .A2(KEYINPUT55), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(KEYINPUT56), .A3(new_n641_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n880_), .B1(new_n889_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n647_), .A2(new_n654_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n552_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n559_), .B1(new_n567_), .B2(new_n555_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n518_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n570_), .B2(new_n518_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n897_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n721_), .B1(new_n896_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n574_), .A2(new_n517_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n644_), .A2(new_n646_), .B1(new_n906_), .B2(new_n900_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n894_), .A2(KEYINPUT56), .A3(new_n641_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n894_), .B2(new_n641_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n756_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT58), .B(new_n907_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n904_), .A2(new_n905_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n721_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n577_), .B(new_n647_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n902_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT57), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n678_), .B1(new_n914_), .B2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT119), .B1(new_n877_), .B2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n901_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n889_), .B2(new_n895_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n713_), .B1(new_n922_), .B2(KEYINPUT58), .ZN(new_n923_));
  INV_X1    g722(.A(new_n913_), .ZN(new_n924_));
  OAI22_X1  g723(.A1(new_n917_), .A2(KEYINPUT57), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n904_), .A2(new_n905_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n679_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n874_), .A2(new_n876_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n920_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n486_), .A2(new_n448_), .A3(new_n509_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(G113gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n934_), .A3(new_n577_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n932_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n938_), .A2(KEYINPUT59), .A3(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n926_), .B1(new_n925_), .B2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n914_), .A2(KEYINPUT121), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n678_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n877_), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n932_), .B(KEYINPUT120), .Z(new_n947_));
  OAI21_X1  g746(.A(new_n941_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n718_), .B1(new_n940_), .B2(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n935_), .B1(new_n949_), .B2(new_n934_), .ZN(G1340gat));
  INV_X1    g749(.A(G120gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n951_), .B1(new_n657_), .B2(KEYINPUT60), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n933_), .B(new_n952_), .C1(KEYINPUT60), .C2(new_n951_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n657_), .B1(new_n940_), .B2(new_n948_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n951_), .ZN(G1341gat));
  INV_X1    g754(.A(G127gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n933_), .A2(new_n956_), .A3(new_n678_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n679_), .B1(new_n940_), .B2(new_n948_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n956_), .ZN(G1342gat));
  INV_X1    g758(.A(G134gat), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n933_), .A2(new_n960_), .A3(new_n915_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n756_), .B1(new_n940_), .B2(new_n948_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n962_), .B2(new_n960_), .ZN(G1343gat));
  NAND3_X1  g762(.A1(new_n454_), .A2(new_n448_), .A3(new_n492_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n486_), .A2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n938_), .A2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n967_), .A2(new_n234_), .A3(new_n577_), .ZN(new_n968_));
  OAI21_X1  g767(.A(G141gat), .B1(new_n966_), .B2(new_n718_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1344gat));
  NAND3_X1  g769(.A1(new_n967_), .A2(new_n235_), .A3(new_n658_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G148gat), .B1(new_n966_), .B2(new_n657_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(G1345gat));
  NAND4_X1  g772(.A1(new_n938_), .A2(KEYINPUT122), .A3(new_n678_), .A4(new_n965_), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n920_), .A2(new_n678_), .A3(new_n930_), .A4(new_n965_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  XNOR2_X1  g776(.A(KEYINPUT61), .B(G155gat), .ZN(new_n978_));
  AND3_X1   g777(.A1(new_n974_), .A2(new_n977_), .A3(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n974_), .B2(new_n977_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1346gat));
  OAI21_X1  g780(.A(G162gat), .B1(new_n966_), .B2(new_n756_), .ZN(new_n982_));
  OR2_X1    g781(.A1(new_n721_), .A2(G162gat), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n982_), .B1(new_n966_), .B2(new_n983_), .ZN(G1347gat));
  NAND3_X1  g783(.A1(new_n486_), .A2(new_n402_), .A3(new_n504_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n985_), .A2(new_n492_), .ZN(new_n986_));
  OAI211_X1 g785(.A(new_n577_), .B(new_n986_), .C1(new_n945_), .C2(new_n877_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n987_), .A2(KEYINPUT123), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n918_), .B1(new_n914_), .B2(KEYINPUT121), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n925_), .A2(new_n942_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n679_), .B1(new_n989_), .B2(new_n990_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n991_), .A2(new_n929_), .ZN(new_n992_));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n993_));
  NAND4_X1  g792(.A1(new_n992_), .A2(new_n993_), .A3(new_n577_), .A4(new_n986_), .ZN(new_n994_));
  NAND3_X1  g793(.A1(new_n988_), .A2(new_n994_), .A3(G169gat), .ZN(new_n995_));
  XNOR2_X1  g794(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n995_), .A2(new_n996_), .ZN(new_n997_));
  INV_X1    g796(.A(new_n996_), .ZN(new_n998_));
  NAND4_X1  g797(.A1(new_n988_), .A2(new_n994_), .A3(G169gat), .A4(new_n998_), .ZN(new_n999_));
  AND2_X1   g798(.A1(new_n992_), .A2(new_n986_), .ZN(new_n1000_));
  NAND4_X1  g799(.A1(new_n1000_), .A2(new_n330_), .A3(new_n332_), .A4(new_n577_), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n997_), .A2(new_n999_), .A3(new_n1001_), .ZN(G1348gat));
  NAND2_X1  g801(.A1(new_n1000_), .A2(new_n658_), .ZN(new_n1003_));
  AND2_X1   g802(.A1(new_n327_), .A2(new_n329_), .ZN(new_n1004_));
  NOR2_X1   g803(.A1(new_n931_), .A2(new_n492_), .ZN(new_n1005_));
  NOR3_X1   g804(.A1(new_n985_), .A2(new_n657_), .A3(new_n309_), .ZN(new_n1006_));
  AOI22_X1  g805(.A1(new_n1003_), .A2(new_n1004_), .B1(new_n1005_), .B2(new_n1006_), .ZN(G1349gat));
  NOR2_X1   g806(.A1(new_n985_), .A2(new_n679_), .ZN(new_n1008_));
  AOI21_X1  g807(.A(G183gat), .B1(new_n1005_), .B2(new_n1008_), .ZN(new_n1009_));
  NOR2_X1   g808(.A1(new_n679_), .A2(new_n352_), .ZN(new_n1010_));
  AOI21_X1  g809(.A(new_n1009_), .B1(new_n1000_), .B2(new_n1010_), .ZN(G1350gat));
  NAND3_X1  g810(.A1(new_n1000_), .A2(new_n353_), .A3(new_n915_), .ZN(new_n1012_));
  AND2_X1   g811(.A1(new_n1000_), .A2(new_n713_), .ZN(new_n1013_));
  OAI21_X1  g812(.A(new_n1012_), .B1(new_n1013_), .B2(new_n303_), .ZN(G1351gat));
  NAND3_X1  g813(.A1(new_n491_), .A2(new_n449_), .A3(new_n504_), .ZN(new_n1015_));
  NOR2_X1   g814(.A1(new_n931_), .A2(new_n1015_), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1016_), .A2(new_n577_), .ZN(new_n1017_));
  XNOR2_X1  g816(.A(new_n1017_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g817(.A1(new_n1016_), .A2(new_n658_), .ZN(new_n1019_));
  XNOR2_X1  g818(.A(new_n1019_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g819(.A(new_n1015_), .ZN(new_n1021_));
  AOI21_X1  g820(.A(new_n679_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1022_));
  XNOR2_X1  g821(.A(new_n1022_), .B(KEYINPUT125), .ZN(new_n1023_));
  NAND4_X1  g822(.A1(new_n920_), .A2(new_n930_), .A3(new_n1021_), .A4(new_n1023_), .ZN(new_n1024_));
  NAND2_X1  g823(.A1(new_n1024_), .A2(KEYINPUT126), .ZN(new_n1025_));
  INV_X1    g824(.A(new_n1025_), .ZN(new_n1026_));
  NOR2_X1   g825(.A1(new_n1024_), .A2(KEYINPUT126), .ZN(new_n1027_));
  OAI22_X1  g826(.A1(new_n1026_), .A2(new_n1027_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1028_));
  INV_X1    g827(.A(new_n1027_), .ZN(new_n1029_));
  NOR2_X1   g828(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1030_));
  NAND3_X1  g829(.A1(new_n1029_), .A2(new_n1030_), .A3(new_n1025_), .ZN(new_n1031_));
  NAND2_X1  g830(.A1(new_n1028_), .A2(new_n1031_), .ZN(G1354gat));
  NAND2_X1  g831(.A1(new_n1016_), .A2(new_n915_), .ZN(new_n1033_));
  XNOR2_X1  g832(.A(KEYINPUT127), .B(G218gat), .ZN(new_n1034_));
  NOR2_X1   g833(.A1(new_n756_), .A2(new_n1034_), .ZN(new_n1035_));
  AOI22_X1  g834(.A1(new_n1033_), .A2(new_n1034_), .B1(new_n1016_), .B2(new_n1035_), .ZN(G1355gat));
endmodule


