//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT72), .ZN(new_n205_));
  INV_X1    g004(.A(G36gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G29gat), .ZN(new_n207_));
  INV_X1    g006(.A(G29gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G36gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT72), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n205_), .A2(new_n210_), .A3(KEYINPUT73), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT73), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(new_n209_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n204_), .A2(KEYINPUT72), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n212_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n203_), .B1(new_n211_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT73), .B1(new_n205_), .B2(new_n210_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n216_), .A3(new_n212_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n202_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(KEYINPUT15), .A3(new_n221_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226_));
  INV_X1    g025(.A(G1gat), .ZN(new_n227_));
  INV_X1    g026(.A(G8gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT14), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G1gat), .B(G8gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n230_), .B(new_n231_), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n224_), .A2(new_n225_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT81), .Z(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(new_n222_), .B2(new_n232_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n222_), .A2(new_n232_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n221_), .A3(new_n218_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n235_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT82), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n234_), .A2(new_n238_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n252_), .A3(new_n248_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n250_), .A2(new_n253_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT83), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(G183gat), .A3(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n255_), .B1(new_n260_), .B2(KEYINPUT23), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(G183gat), .B2(G190gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT84), .B(G176gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT22), .B(G169gat), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n263_), .A2(new_n264_), .B1(G169gat), .B2(G176gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT25), .B(G183gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(G190gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(G169gat), .B2(G176gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(G169gat), .B2(G176gat), .ZN(new_n273_));
  INV_X1    g072(.A(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(G176gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n270_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT23), .B1(new_n257_), .B2(new_n259_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n256_), .A2(KEYINPUT23), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n262_), .A2(new_n265_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282_));
  INV_X1    g081(.A(G43gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G127gat), .B(G134gat), .Z(new_n286_));
  XOR2_X1   g085(.A(G113gat), .B(G120gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n285_), .B(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G227gat), .A2(G233gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(G15gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT30), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT31), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n294_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G197gat), .A2(G204gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G197gat), .A2(G204gat), .ZN(new_n301_));
  OR3_X1    g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT90), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT90), .B1(new_n300_), .B2(new_n301_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G211gat), .B(G218gat), .Z(new_n304_));
  NAND4_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT21), .A4(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(G197gat), .A2(G204gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(KEYINPUT21), .A3(new_n299_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n306_), .A2(KEYINPUT88), .A3(KEYINPUT21), .A4(new_n299_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT21), .B1(new_n306_), .B2(new_n299_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(new_n304_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n305_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n322_), .A2(new_n325_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G155gat), .ZN(new_n331_));
  INV_X1    g130(.A(G162gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT85), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(G155gat), .B2(G162gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n330_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n328_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G141gat), .B(G148gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(KEYINPUT1), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(G155gat), .A3(G162gat), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(new_n335_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n338_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n317_), .B1(new_n318_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(G228gat), .A3(G233gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT86), .B1(new_n337_), .B2(new_n344_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n338_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n333_), .A2(new_n335_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n339_), .A2(new_n341_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n328_), .A2(new_n336_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n349_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n317_), .B(new_n348_), .C1(new_n318_), .C2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n347_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT91), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n347_), .A2(new_n363_), .A3(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n357_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n367_));
  OR3_X1    g166(.A1(new_n366_), .A2(KEYINPUT29), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n366_), .B2(KEYINPUT29), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G22gat), .B(G50gat), .Z(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n368_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n365_), .A2(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n362_), .A2(new_n372_), .A3(new_n374_), .A4(new_n364_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n286_), .B(new_n287_), .Z(new_n379_));
  NAND3_X1  g178(.A1(new_n349_), .A2(new_n379_), .A3(new_n356_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n345_), .A2(new_n288_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT95), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n380_), .A2(KEYINPUT95), .A3(new_n381_), .A4(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n380_), .A2(KEYINPUT4), .A3(new_n382_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n349_), .A2(new_n356_), .A3(new_n379_), .A4(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n388_), .A2(G225gat), .A3(G233gat), .A4(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G57gat), .B(G85gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT94), .ZN(new_n394_));
  XOR2_X1   g193(.A(G1gat), .B(G29gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n392_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n387_), .A2(new_n398_), .A3(new_n391_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT19), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n262_), .A2(new_n265_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n277_), .A2(new_n280_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n408_), .ZN(new_n409_));
  OAI22_X1  g208(.A1(new_n278_), .A2(new_n279_), .B1(G183gat), .B2(G190gat), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n277_), .A2(new_n261_), .B1(new_n265_), .B2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n300_), .A2(new_n301_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT88), .B1(new_n412_), .B2(KEYINPUT21), .ZN(new_n413_));
  INV_X1    g212(.A(new_n310_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n314_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT89), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n411_), .B1(new_n418_), .B2(new_n305_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n405_), .B1(new_n409_), .B2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G8gat), .B(G36gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n427_));
  INV_X1    g226(.A(new_n305_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n411_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n317_), .A2(new_n408_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n405_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(KEYINPUT20), .A4(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n420_), .A2(new_n427_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n411_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n281_), .B1(new_n418_), .B2(new_n305_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n405_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n429_), .B2(new_n281_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n317_), .A2(new_n435_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n432_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n427_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n434_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n392_), .A2(KEYINPUT97), .A3(new_n399_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n403_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n402_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n387_), .A2(KEYINPUT33), .A3(new_n391_), .A4(new_n398_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n436_), .A2(new_n437_), .A3(new_n405_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n432_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n425_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n380_), .A2(new_n382_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n381_), .B1(new_n454_), .B2(KEYINPUT96), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(KEYINPUT96), .B2(new_n454_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n388_), .A2(new_n381_), .A3(new_n390_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n399_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n420_), .A2(new_n426_), .A3(new_n433_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n450_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n378_), .B1(new_n446_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n402_), .A2(new_n401_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n398_), .B1(new_n387_), .B2(new_n391_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n445_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n463_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n459_), .A2(KEYINPUT27), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n426_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT27), .B1(new_n453_), .B2(new_n459_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n376_), .A2(new_n377_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n403_), .A2(KEYINPUT98), .A3(new_n445_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n468_), .A2(new_n473_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n298_), .B1(new_n462_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n468_), .A2(new_n475_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n378_), .A2(new_n298_), .A3(new_n473_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n477_), .A2(KEYINPUT99), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n462_), .A2(new_n476_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n297_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT99), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n254_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G71gat), .B(G78gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT11), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n490_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT66), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n497_), .B(new_n490_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n505_), .B(KEYINPUT7), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n508_), .B(KEYINPUT6), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(KEYINPUT65), .A3(new_n504_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n513_), .A2(KEYINPUT8), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT10), .B(G99gat), .Z(new_n520_));
  AOI21_X1  g319(.A(new_n510_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n503_), .A2(KEYINPUT64), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT64), .B1(new_n503_), .B2(new_n522_), .ZN(new_n524_));
  OAI221_X1 g323(.A(new_n502_), .B1(new_n522_), .B2(new_n503_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n513_), .B2(KEYINPUT8), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n499_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT65), .B1(new_n516_), .B2(new_n504_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT8), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n530_), .A2(new_n531_), .B1(new_n525_), .B2(new_n521_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n513_), .A2(new_n517_), .A3(KEYINPUT8), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(KEYINPUT12), .B(new_n490_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n528_), .A2(new_n529_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n532_), .A2(new_n533_), .A3(new_n498_), .A4(new_n496_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT68), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n528_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n540_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n545_), .B(new_n546_), .C1(new_n544_), .C2(new_n538_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G120gat), .B(G148gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n543_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n543_), .A2(new_n547_), .A3(KEYINPUT70), .A4(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n551_), .B(KEYINPUT69), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT13), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n562_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT34), .Z(new_n568_));
  INV_X1    g367(.A(KEYINPUT35), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n222_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT74), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n569_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n224_), .A2(new_n534_), .A3(new_n225_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n572_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n570_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT75), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n570_), .B(KEYINPUT76), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n575_), .A2(new_n573_), .A3(new_n571_), .A4(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n578_), .A2(new_n579_), .A3(new_n583_), .A4(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT78), .ZN(new_n587_));
  INV_X1    g386(.A(new_n585_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n577_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n590_), .B2(new_n570_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n583_), .B(KEYINPUT36), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT77), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n586_), .B(new_n587_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT79), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n232_), .B(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(new_n495_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(new_n495_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n600_), .A2(KEYINPUT17), .A3(new_n605_), .A4(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n605_), .B(KEYINPUT17), .Z(new_n608_));
  OR2_X1    g407(.A1(new_n599_), .A2(new_n499_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n599_), .A2(new_n499_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n578_), .A2(new_n585_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n593_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n616_), .A2(new_n587_), .A3(KEYINPUT37), .A4(new_n586_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n596_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n487_), .A2(new_n566_), .A3(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n620_), .A2(G1gat), .A3(new_n479_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n616_), .A2(new_n586_), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n612_), .B(new_n624_), .C1(new_n482_), .C2(new_n486_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n563_), .A2(new_n565_), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n558_), .B(new_n560_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(new_n254_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n479_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n622_), .A2(new_n623_), .A3(new_n631_), .ZN(G1324gat));
  NOR3_X1   g431(.A1(new_n620_), .A2(G8gat), .A3(new_n473_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G8gat), .B1(new_n630_), .B2(new_n473_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT39), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n636_), .B(G8gat), .C1(new_n630_), .C2(new_n473_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n638_), .B(new_n640_), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n630_), .B2(new_n297_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT41), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n620_), .A2(G15gat), .A3(new_n297_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  OR3_X1    g444(.A1(new_n620_), .A2(G22gat), .A3(new_n378_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n625_), .A2(new_n474_), .A3(new_n629_), .ZN(new_n647_));
  XOR2_X1   g446(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(G22gat), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G22gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n624_), .A2(new_n612_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT103), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n628_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n487_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n478_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n596_), .A2(new_n617_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n483_), .A2(KEYINPUT99), .A3(new_n297_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n481_), .A2(new_n479_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n477_), .A2(KEYINPUT99), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT43), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n482_), .A2(new_n486_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n658_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n254_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n566_), .A2(new_n669_), .A3(new_n612_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT102), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n674_), .B(new_n671_), .C1(new_n664_), .C2(new_n667_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n479_), .A2(new_n208_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n657_), .B1(new_n676_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  INV_X1    g478(.A(new_n473_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n206_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n473_), .A2(G36gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT104), .B1(new_n655_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n487_), .A2(new_n685_), .A3(new_n654_), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n679_), .B1(new_n681_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n687_), .B(KEYINPUT45), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n673_), .A2(new_n675_), .A3(new_n473_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n691_), .B(KEYINPUT46), .C1(new_n206_), .C2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1329gat));
  INV_X1    g493(.A(new_n673_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n672_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n695_), .A2(G43gat), .A3(new_n298_), .A4(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n283_), .B1(new_n655_), .B2(new_n297_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT47), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n701_), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n676_), .B2(new_n474_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n655_), .A2(G50gat), .A3(new_n378_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT105), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708_));
  INV_X1    g507(.A(new_n706_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n673_), .A2(new_n675_), .A3(new_n378_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n708_), .B(new_n709_), .C1(new_n710_), .C2(new_n704_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(G1331gat));
  NAND3_X1  g511(.A1(new_n625_), .A2(new_n254_), .A3(new_n628_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n479_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n669_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n566_), .A2(new_n618_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n479_), .A2(G57gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1332gat));
  OR3_X1    g518(.A1(new_n717_), .A2(G64gat), .A3(new_n473_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G64gat), .B1(new_n713_), .B2(new_n473_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT48), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT48), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT106), .B(new_n720_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1333gat));
  NOR2_X1   g527(.A1(new_n297_), .A2(G71gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT107), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n715_), .A2(new_n716_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G71gat), .B1(new_n713_), .B2(new_n297_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(KEYINPUT49), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(KEYINPUT49), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT108), .B(new_n731_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n713_), .B2(new_n378_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n378_), .A2(G78gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n717_), .B2(new_n742_), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n653_), .A2(new_n566_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n715_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n500_), .A3(new_n478_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n566_), .A2(new_n669_), .A3(new_n613_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n666_), .B1(new_n665_), .B2(new_n658_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n596_), .A2(new_n617_), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT43), .B(new_n750_), .C1(new_n482_), .C2(new_n486_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n668_), .A2(KEYINPUT109), .A3(new_n748_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n479_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n747_), .B1(new_n756_), .B2(new_n500_), .ZN(G1336gat));
  OAI21_X1  g556(.A(new_n501_), .B1(new_n745_), .B2(new_n473_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT110), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n754_), .A2(new_n755_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n473_), .A2(new_n501_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(G1337gat));
  INV_X1    g561(.A(G99gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n760_), .B2(new_n298_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n298_), .A2(new_n520_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n745_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT51), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n297_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n769_));
  OAI221_X1 g568(.A(new_n768_), .B1(new_n745_), .B2(new_n765_), .C1(new_n769_), .C2(new_n763_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n746_), .A2(new_n519_), .A3(new_n474_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n668_), .A2(new_n474_), .A3(new_n748_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G106gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n772_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  AOI21_X1  g580(.A(new_n254_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n543_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n536_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n532_), .A2(new_n533_), .B1(new_n498_), .B2(new_n496_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n785_), .B(new_n538_), .C1(new_n786_), .C2(KEYINPUT12), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n528_), .A2(new_n529_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(KEYINPUT113), .A3(new_n785_), .A4(new_n538_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n791_), .A3(new_n546_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT55), .B(new_n537_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n784_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n557_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n795_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n782_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n563_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n237_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n248_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n234_), .A2(new_n240_), .A3(new_n237_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n801_), .B2(new_n248_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n252_), .B1(new_n251_), .B2(new_n248_), .ZN(new_n807_));
  AND4_X1   g606(.A1(new_n252_), .A2(new_n239_), .A3(new_n244_), .A4(new_n248_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n806_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n800_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n624_), .B1(new_n799_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n809_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n815_), .B(new_n817_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n658_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n794_), .A2(new_n795_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n796_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n817_), .B1(new_n823_), .B2(new_n815_), .ZN(new_n824_));
  OAI22_X1  g623(.A1(new_n812_), .A2(new_n814_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n823_), .A2(new_n782_), .B1(new_n800_), .B2(new_n810_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n826_), .A2(new_n624_), .A3(new_n813_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n612_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n750_), .A2(new_n566_), .A3(new_n254_), .A4(new_n613_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n619_), .A2(new_n566_), .A3(new_n254_), .A4(new_n831_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(KEYINPUT112), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT112), .B1(new_n834_), .B2(new_n835_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n828_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n479_), .A2(new_n480_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n838_), .A2(new_n839_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n839_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n838_), .A2(KEYINPUT117), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n828_), .B(new_n848_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n841_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n845_), .B(new_n669_), .C1(new_n846_), .C2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G113gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n840_), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n854_), .A2(G113gat), .A3(new_n254_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(G1340gat));
  OAI211_X1 g655(.A(new_n845_), .B(new_n628_), .C1(new_n846_), .C2(new_n850_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G120gat), .ZN(new_n858_));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n566_), .B2(KEYINPUT60), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(KEYINPUT60), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(KEYINPUT119), .B2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n850_), .B(new_n862_), .C1(KEYINPUT119), .C2(new_n860_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n863_), .ZN(G1341gat));
  OAI211_X1 g663(.A(new_n845_), .B(new_n613_), .C1(new_n846_), .C2(new_n850_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G127gat), .ZN(new_n866_));
  OR3_X1    g665(.A1(new_n854_), .A2(G127gat), .A3(new_n612_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1342gat));
  INV_X1    g667(.A(new_n624_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n869_), .B(new_n841_), .C1(new_n847_), .C2(new_n849_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n870_), .B2(G134gat), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  INV_X1    g671(.A(G134gat), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n872_), .B(new_n873_), .C1(new_n854_), .C2(new_n869_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n834_), .A2(new_n835_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n834_), .A2(KEYINPUT112), .A3(new_n835_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n813_), .B1(new_n826_), .B2(new_n624_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n812_), .A2(new_n814_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n879_), .B(new_n880_), .C1(new_n824_), .C2(new_n819_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n877_), .A2(new_n878_), .B1(new_n881_), .B2(new_n612_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n842_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT118), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n838_), .A2(new_n839_), .A3(new_n842_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n854_), .B2(KEYINPUT59), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT121), .B(G134gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n750_), .A2(new_n888_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n871_), .A2(new_n874_), .B1(new_n887_), .B2(new_n889_), .ZN(G1343gat));
  NOR3_X1   g689(.A1(new_n680_), .A2(new_n378_), .A3(new_n298_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n478_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n669_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n628_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g696(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n892_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n877_), .A2(new_n878_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n848_), .B1(new_n901_), .B2(new_n828_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n849_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n613_), .B(new_n900_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT61), .B(G155gat), .Z(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n905_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n893_), .B2(new_n613_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n899_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(new_n905_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n893_), .A2(new_n613_), .A3(new_n907_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n898_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(G1346gat));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914_));
  AOI21_X1  g713(.A(G162gat), .B1(new_n893_), .B2(new_n624_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n658_), .A2(G162gat), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(KEYINPUT124), .Z(new_n917_));
  AND3_X1   g716(.A1(new_n853_), .A2(new_n900_), .A3(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n914_), .B1(new_n915_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n893_), .A2(new_n917_), .ZN(new_n920_));
  AOI211_X1 g719(.A(new_n869_), .B(new_n892_), .C1(new_n847_), .C2(new_n849_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n920_), .B(KEYINPUT125), .C1(new_n921_), .C2(G162gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n922_), .ZN(G1347gat));
  NOR4_X1   g722(.A1(new_n478_), .A2(new_n297_), .A3(new_n474_), .A4(new_n473_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n838_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n274_), .B1(new_n926_), .B2(new_n669_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n927_), .A2(KEYINPUT62), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n669_), .A3(new_n264_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(KEYINPUT62), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(new_n929_), .A3(new_n930_), .ZN(G1348gat));
  NAND4_X1  g730(.A1(new_n853_), .A2(G176gat), .A3(new_n628_), .A4(new_n924_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT126), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n263_), .B1(new_n925_), .B2(new_n566_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n932_), .A2(KEYINPUT126), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1349gat));
  NOR3_X1   g736(.A1(new_n925_), .A2(new_n266_), .A3(new_n612_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n853_), .A2(new_n613_), .A3(new_n924_), .ZN(new_n939_));
  INV_X1    g738(.A(G183gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n925_), .B2(new_n750_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n624_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n925_), .B2(new_n943_), .ZN(G1351gat));
  NOR4_X1   g743(.A1(new_n478_), .A2(new_n378_), .A3(new_n298_), .A4(new_n473_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n669_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n628_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g750(.A(new_n612_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n947_), .A2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(KEYINPUT127), .ZN(new_n955_));
  XOR2_X1   g754(.A(new_n953_), .B(new_n955_), .Z(G1354gat));
  INV_X1    g755(.A(new_n947_), .ZN(new_n957_));
  OR3_X1    g756(.A1(new_n957_), .A2(G218gat), .A3(new_n869_), .ZN(new_n958_));
  OAI21_X1  g757(.A(G218gat), .B1(new_n957_), .B2(new_n750_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1355gat));
endmodule


