//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(KEYINPUT81), .A3(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n204_), .B1(KEYINPUT81), .B2(G169gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n203_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n211_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT23), .A3(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT82), .A4(new_n213_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n209_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT25), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT78), .A3(G183gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n232_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT24), .A3(new_n203_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n231_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n218_), .A2(new_n219_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n210_), .A2(new_n213_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n238_), .A2(new_n239_), .B1(new_n240_), .B2(new_n211_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n202_), .B1(new_n225_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n238_), .ZN(new_n244_));
  AND2_X1   g043(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n245_));
  NOR2_X1   g044(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n244_), .B1(new_n212_), .B2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n236_), .A2(new_n234_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n231_), .A3(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n221_), .A2(new_n220_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n223_), .B1(new_n251_), .B2(new_n216_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(KEYINPUT83), .C1(new_n252_), .C2(new_n209_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n243_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G71gat), .B(G99gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT85), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G15gat), .B(G43gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n254_), .B(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G127gat), .B(G134gat), .Z(new_n260_));
  XOR2_X1   g059(.A(G113gat), .B(G120gat), .Z(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT86), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G113gat), .B(G120gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(KEYINPUT86), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n259_), .B(new_n269_), .Z(new_n270_));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT84), .Z(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT30), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT31), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n270_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G22gat), .B(G50gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n276_), .B(KEYINPUT93), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(KEYINPUT88), .A2(G141gat), .A3(G148gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT2), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n284_), .A2(new_n285_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n283_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n287_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n279_), .B2(KEYINPUT1), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n279_), .A2(new_n299_), .A3(KEYINPUT1), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n281_), .B1(new_n280_), .B2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n298_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT29), .B1(new_n294_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT21), .B1(new_n308_), .B2(KEYINPUT92), .ZN(new_n309_));
  INV_X1    g108(.A(G218gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G211gat), .ZN(new_n311_));
  INV_X1    g110(.A(G211gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G218gat), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n311_), .A2(new_n313_), .A3(KEYINPUT92), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G197gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT90), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G197gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n319_), .A3(G204gat), .ZN(new_n320_));
  INV_X1    g119(.A(G204gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n316_), .B2(G204gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n315_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n311_), .A2(new_n313_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(G197gat), .B2(G204gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n320_), .A2(new_n329_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G106gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n307_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  OR2_X1    g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT3), .B1(new_n338_), .B2(KEYINPUT88), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n339_), .A2(new_n293_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n282_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n302_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n305_), .B1(new_n342_), .B2(new_n300_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n297_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n337_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n315_), .A2(new_n325_), .B1(new_n332_), .B2(new_n331_), .ZN(new_n346_));
  OAI21_X1  g145(.A(G106gat), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(G78gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n336_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n336_), .B2(new_n347_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n340_), .A2(new_n282_), .B1(new_n343_), .B2(new_n297_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n337_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n355_), .B(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n352_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n355_), .B(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n336_), .A2(new_n347_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n350_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(new_n351_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n278_), .B1(new_n359_), .B2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n358_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n351_), .A3(new_n360_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n277_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n344_), .A2(new_n341_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n262_), .A2(new_n266_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n341_), .A2(new_n344_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT4), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n269_), .B1(new_n306_), .B2(new_n294_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G85gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT0), .B(G57gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n354_), .A2(new_n372_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n377_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n375_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n380_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n384_), .B1(new_n380_), .B2(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT100), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AND4_X1   g190(.A1(new_n390_), .A2(new_n380_), .A3(new_n384_), .A4(new_n387_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n221_), .A2(new_n220_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT82), .B1(new_n247_), .B2(new_n212_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n233_), .A2(KEYINPUT94), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT94), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT24), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n203_), .A3(new_n235_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT25), .B(G183gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n226_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n397_), .A2(new_n399_), .A3(new_n232_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT95), .B1(new_n396_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n235_), .A2(new_n203_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n404_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n222_), .A2(new_n410_), .A3(new_n411_), .A4(new_n403_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n206_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n203_), .B(new_n414_), .C1(new_n241_), .C2(new_n223_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n406_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n334_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT96), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n243_), .A2(new_n253_), .A3(new_n346_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n420_), .A3(new_n334_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n418_), .A2(KEYINPUT20), .A3(new_n419_), .A4(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT19), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT20), .B(new_n426_), .C1(new_n416_), .C2(new_n334_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n346_), .B1(new_n243_), .B2(new_n253_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT18), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n432_), .B(new_n433_), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT99), .B(KEYINPUT20), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n346_), .A2(new_n415_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n396_), .A2(new_n405_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n424_), .B1(new_n428_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT32), .A3(new_n434_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n393_), .A2(new_n436_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n386_), .A2(KEYINPUT97), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT97), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n377_), .A2(new_n385_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n376_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n384_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT98), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT98), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n452_), .A3(new_n384_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n374_), .A2(new_n379_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n451_), .B(new_n453_), .C1(new_n376_), .C2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n389_), .B(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n425_), .A2(new_n434_), .A3(new_n430_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n434_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n416_), .A2(new_n420_), .A3(new_n334_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n420_), .B1(new_n416_), .B2(new_n334_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n419_), .A2(KEYINPUT20), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n426_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n459_), .B1(new_n464_), .B2(new_n429_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .A4(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n370_), .B1(new_n445_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n458_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n365_), .B(new_n368_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n419_), .A2(KEYINPUT20), .ZN(new_n474_));
  NOR4_X1   g273(.A1(new_n474_), .A2(new_n460_), .A3(new_n461_), .A4(new_n424_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n442_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n459_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  AND4_X1   g276(.A1(KEYINPUT101), .A2(new_n477_), .A3(KEYINPUT27), .A4(new_n458_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT27), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n443_), .B2(new_n459_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT101), .B1(new_n480_), .B2(new_n458_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n471_), .B(new_n473_), .C1(new_n478_), .C2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n467_), .B1(new_n482_), .B2(KEYINPUT103), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n469_), .B1(new_n465_), .B2(new_n458_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(new_n472_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT103), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n485_), .B(new_n486_), .C1(new_n481_), .C2(new_n478_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n275_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n393_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n275_), .A2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n471_), .B(new_n369_), .C1(new_n478_), .C2(new_n481_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n494_));
  XOR2_X1   g293(.A(G120gat), .B(G148gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(G176gat), .B(G204gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n501_), .A2(new_n502_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT12), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT6), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  INV_X1    g317(.A(G99gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n335_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n512_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT8), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT65), .B1(new_n514_), .B2(new_n516_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n514_), .A2(new_n516_), .A3(KEYINPUT65), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n522_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n512_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n524_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n527_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n511_), .B1(new_n510_), .B2(KEYINPUT9), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT64), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n533_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT10), .B(G99gat), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n335_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n531_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n508_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n505_), .A2(new_n506_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n522_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n527_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(new_n525_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n530_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n547_), .A2(new_n548_), .B1(new_n523_), .B2(KEYINPUT8), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n532_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT66), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n531_), .A2(new_n552_), .A3(new_n541_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n544_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n543_), .B1(new_n554_), .B2(KEYINPUT12), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n551_), .A2(new_n553_), .A3(new_n544_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(KEYINPUT67), .A3(new_n557_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n555_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n544_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT66), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n552_), .B1(new_n531_), .B2(new_n541_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n557_), .B1(new_n566_), .B2(new_n556_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n499_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT12), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n566_), .A2(new_n569_), .B1(new_n542_), .B2(new_n508_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n561_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT67), .B1(new_n556_), .B2(new_n557_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n567_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n499_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT69), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n568_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(KEYINPUT69), .B(new_n499_), .C1(new_n562_), .C2(new_n567_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT13), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT13), .B1(new_n578_), .B2(new_n579_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n494_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n579_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT13), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT70), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G15gat), .B(G22gat), .ZN(new_n589_));
  INV_X1    g388(.A(G1gat), .ZN(new_n590_));
  INV_X1    g389(.A(G8gat), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT14), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G1gat), .B(G8gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G29gat), .B(G36gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G43gat), .B(G50gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n595_), .B(new_n598_), .Z(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n598_), .B(KEYINPUT15), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n595_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n595_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n598_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n606_), .A3(new_n600_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G169gat), .B(G197gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n602_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(KEYINPUT76), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT76), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n616_), .A3(new_n612_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT77), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT34), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT35), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT72), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(KEYINPUT35), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n625_), .B(new_n626_), .C1(new_n542_), .C2(new_n603_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n551_), .A2(new_n553_), .A3(new_n598_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n624_), .A3(new_n623_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n624_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n631_), .A3(new_n628_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT36), .Z(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT73), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n632_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT74), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n630_), .A2(new_n632_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n635_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n638_), .A2(KEYINPUT74), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT37), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n630_), .A2(new_n636_), .A3(new_n632_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n595_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(new_n563_), .ZN(new_n653_));
  XOR2_X1   g452(.A(G127gat), .B(G155gat), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT16), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G183gat), .B(G211gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT17), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n653_), .A2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT75), .Z(new_n661_));
  AND2_X1   g460(.A1(new_n657_), .A2(new_n658_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n653_), .A2(new_n659_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n650_), .A2(new_n665_), .ZN(new_n666_));
  NOR4_X1   g465(.A1(new_n493_), .A2(new_n588_), .A3(new_n620_), .A4(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n590_), .A3(new_n393_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n478_), .A2(new_n481_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n473_), .A2(new_n471_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT103), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n467_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n487_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n275_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n492_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n618_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n588_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n677_), .A2(new_n648_), .A3(new_n665_), .A4(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n680_), .B2(new_n489_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n668_), .A2(new_n681_), .ZN(new_n682_));
  MUX2_X1   g481(.A(new_n668_), .B(new_n682_), .S(KEYINPUT38), .Z(G1324gat));
  NOR2_X1   g482(.A1(new_n669_), .A2(new_n484_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G8gat), .B1(new_n680_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT39), .ZN(new_n686_));
  INV_X1    g485(.A(new_n684_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n667_), .A2(new_n591_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n689_), .B(new_n691_), .ZN(G1325gat));
  OAI21_X1  g491(.A(G15gat), .B1(new_n680_), .B2(new_n674_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT41), .Z(new_n694_));
  INV_X1    g493(.A(G15gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n667_), .A2(new_n695_), .A3(new_n275_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1326gat));
  OAI21_X1  g496(.A(G22gat), .B1(new_n680_), .B2(new_n369_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT42), .ZN(new_n699_));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n667_), .A2(new_n700_), .A3(new_n370_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1327gat));
  NOR2_X1   g501(.A1(new_n665_), .A2(new_n648_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n582_), .A2(new_n587_), .A3(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n704_), .B(new_n619_), .C1(new_n488_), .C2(new_n492_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n677_), .A2(KEYINPUT106), .A3(new_n619_), .A4(new_n704_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n393_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n650_), .B(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n650_), .A2(KEYINPUT43), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n714_), .A2(KEYINPUT43), .B1(new_n677_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n679_), .A2(new_n664_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n711_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n717_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n677_), .B2(new_n713_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n715_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n493_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n719_), .C1(new_n721_), .C2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n718_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n393_), .A2(G29gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n710_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT107), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT107), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n718_), .A2(new_n687_), .A3(new_n724_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G36gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n684_), .A2(G36gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n707_), .A2(new_n708_), .A3(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT45), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n729_), .B(new_n730_), .C1(new_n732_), .C2(new_n735_), .ZN(new_n736_));
  AND4_X1   g535(.A1(KEYINPUT107), .A2(new_n732_), .A3(new_n728_), .A4(new_n735_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n718_), .A2(G43gat), .A3(new_n724_), .A4(new_n275_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n707_), .A2(new_n708_), .A3(new_n275_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741_));
  INV_X1    g540(.A(G43gat), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n739_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g545(.A1(new_n369_), .A2(G50gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT110), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n709_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n725_), .A2(KEYINPUT109), .A3(new_n370_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT109), .B1(new_n725_), .B2(new_n370_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n751_), .B2(new_n752_), .ZN(G1331gat));
  NAND2_X1  g552(.A1(new_n677_), .A2(new_n678_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n582_), .A2(new_n587_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n664_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n650_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n754_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT111), .ZN(new_n759_));
  INV_X1    g558(.A(G57gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n393_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n648_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n493_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n620_), .A4(new_n756_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n677_), .A2(new_n648_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n756_), .A2(new_n620_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT112), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n765_), .A2(new_n768_), .A3(new_n393_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n760_), .B2(new_n769_), .ZN(G1332gat));
  INV_X1    g569(.A(G64gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n759_), .A2(new_n771_), .A3(new_n687_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n765_), .A2(new_n768_), .A3(new_n687_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G64gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G64gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1333gat));
  NOR2_X1   g576(.A1(new_n674_), .A2(G71gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n759_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n768_), .A3(new_n275_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G71gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G71gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT113), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n779_), .B(new_n786_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1334gat));
  NAND3_X1  g587(.A1(new_n759_), .A2(new_n349_), .A3(new_n370_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n765_), .A2(new_n768_), .A3(new_n370_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G78gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G78gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(G1335gat));
  NOR2_X1   g593(.A1(new_n665_), .A2(new_n618_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n588_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT114), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n716_), .A2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT115), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n393_), .A2(G85gat), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT116), .Z(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n677_), .A2(new_n678_), .A3(new_n588_), .A4(new_n703_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n393_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n802_), .A2(new_n805_), .ZN(G1336gat));
  OAI21_X1  g605(.A(G92gat), .B1(new_n799_), .B2(new_n684_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n803_), .A2(G92gat), .A3(new_n684_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1337gat));
  NOR3_X1   g608(.A1(new_n716_), .A2(new_n797_), .A3(new_n674_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n275_), .A2(new_n539_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n810_), .A2(new_n519_), .B1(new_n803_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n804_), .A2(new_n335_), .A3(new_n370_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815_));
  INV_X1    g614(.A(new_n797_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n370_), .C1(new_n721_), .C2(new_n723_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n817_), .B2(G106gat), .ZN(new_n818_));
  AOI211_X1 g617(.A(KEYINPUT52), .B(new_n335_), .C1(new_n798_), .C2(new_n370_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n814_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT53), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n814_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n666_), .A2(new_n619_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n585_), .A2(new_n586_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n599_), .A2(new_n600_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n604_), .A2(new_n606_), .A3(new_n601_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n612_), .ZN(new_n835_));
  AND4_X1   g634(.A1(new_n614_), .A2(new_n578_), .A3(new_n579_), .A4(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT117), .B1(new_n618_), .B2(new_n576_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n618_), .A2(KEYINPUT117), .A3(new_n576_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n556_), .B(new_n543_), .C1(new_n554_), .C2(KEYINPUT12), .ZN(new_n840_));
  INV_X1    g639(.A(new_n557_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n562_), .B2(KEYINPUT55), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n570_), .B(KEYINPUT55), .C1(new_n571_), .C2(new_n572_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n499_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT118), .B1(new_n847_), .B2(KEYINPUT119), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n838_), .A2(new_n839_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT118), .B(new_n499_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n836_), .B1(new_n849_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n832_), .B1(new_n854_), .B2(new_n762_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n839_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n573_), .A2(new_n857_), .B1(new_n841_), .B2(new_n840_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n575_), .B1(new_n858_), .B2(new_n844_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n848_), .ZN(new_n860_));
  OAI22_X1  g659(.A1(new_n856_), .A2(new_n837_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n852_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n648_), .C1(new_n862_), .C2(new_n836_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n576_), .A2(new_n614_), .A3(new_n835_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n865_));
  NOR2_X1   g664(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n859_), .B2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n846_), .A2(new_n866_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n650_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT58), .B(new_n864_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n855_), .A2(new_n863_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n664_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n876_), .A2(KEYINPUT121), .A3(new_n664_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n831_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n674_), .A2(new_n489_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n491_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(KEYINPUT59), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n825_), .B1(new_n881_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n831_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n877_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n884_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT59), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n876_), .A2(KEYINPUT121), .A3(new_n664_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT121), .B1(new_n876_), .B2(new_n664_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n888_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(KEYINPUT122), .A3(new_n885_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n887_), .A2(new_n619_), .A3(new_n892_), .A4(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G113gat), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n891_), .A2(G113gat), .A3(new_n678_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1340gat));
  NAND4_X1  g699(.A1(new_n887_), .A2(new_n588_), .A3(new_n892_), .A4(new_n896_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G120gat), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n755_), .A2(KEYINPUT60), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n903_), .B(KEYINPUT60), .S(G120gat), .Z(new_n904_));
  NAND3_X1  g703(.A1(new_n889_), .A2(new_n890_), .A3(new_n904_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT123), .Z(new_n906_));
  NAND2_X1  g705(.A1(new_n902_), .A2(new_n906_), .ZN(G1341gat));
  NAND4_X1  g706(.A1(new_n887_), .A2(new_n665_), .A3(new_n892_), .A4(new_n896_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G127gat), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n891_), .A2(G127gat), .A3(new_n664_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1342gat));
  NAND4_X1  g710(.A1(new_n887_), .A2(new_n873_), .A3(new_n892_), .A4(new_n896_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G134gat), .ZN(new_n913_));
  OR3_X1    g712(.A1(new_n891_), .A2(G134gat), .A3(new_n648_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1343gat));
  NOR3_X1   g714(.A1(new_n275_), .A2(new_n489_), .A3(new_n369_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n684_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n888_), .B2(new_n877_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n618_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n588_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n665_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT124), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n918_), .A2(new_n925_), .A3(new_n665_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT61), .B(G155gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  AOI21_X1  g728(.A(G162gat), .B1(new_n918_), .B2(new_n762_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n713_), .A2(G162gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n918_), .B2(new_n931_), .ZN(G1347gat));
  NOR3_X1   g731(.A1(new_n684_), .A2(new_n490_), .A3(new_n370_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n895_), .A2(new_n618_), .A3(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G169gat), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n895_), .A2(new_n933_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n938_), .A2(new_n413_), .A3(new_n618_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n934_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n937_), .A2(new_n939_), .A3(new_n940_), .ZN(G1348gat));
  NAND4_X1  g740(.A1(new_n889_), .A2(G176gat), .A3(new_n588_), .A4(new_n933_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT126), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n895_), .A2(new_n588_), .A3(new_n933_), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n944_), .A2(KEYINPUT125), .A3(new_n206_), .ZN(new_n945_));
  AOI21_X1  g744(.A(KEYINPUT125), .B1(new_n944_), .B2(new_n206_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n943_), .A2(new_n945_), .A3(new_n946_), .ZN(G1349gat));
  AND2_X1   g746(.A1(new_n889_), .A2(new_n933_), .ZN(new_n948_));
  AOI21_X1  g747(.A(G183gat), .B1(new_n948_), .B2(new_n665_), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n664_), .A2(new_n402_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n938_), .B2(new_n951_), .ZN(G1350gat));
  NAND2_X1  g751(.A1(new_n938_), .A2(new_n873_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(G190gat), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n938_), .A2(new_n226_), .A3(new_n762_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n684_), .A2(new_n275_), .A3(new_n472_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n889_), .A2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n618_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n588_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g761(.A1(new_n958_), .A2(new_n665_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  AND2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n963_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n966_), .B1(new_n963_), .B2(new_n964_), .ZN(G1354gat));
  NAND2_X1  g766(.A1(new_n958_), .A2(new_n762_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(KEYINPUT127), .B(G218gat), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n650_), .A2(new_n969_), .ZN(new_n970_));
  AOI22_X1  g769(.A1(new_n968_), .A2(new_n969_), .B1(new_n958_), .B2(new_n970_), .ZN(G1355gat));
endmodule


