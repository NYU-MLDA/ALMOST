//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  AND2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT86), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G155gat), .ZN(new_n211_));
  INV_X1    g010(.A(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT86), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n218_), .A2(new_n221_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  INV_X1    g025(.A(G141gat), .ZN(new_n227_));
  INV_X1    g026(.A(G148gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT3), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n224_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n217_), .B1(new_n223_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n228_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n233_));
  AND4_X1   g032(.A1(new_n220_), .A2(new_n232_), .A3(new_n222_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n213_), .A2(new_n235_), .A3(new_n215_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n207_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n210_), .A2(new_n216_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n229_), .A2(new_n226_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n224_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n223_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n205_), .B(new_n206_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n234_), .A2(new_n236_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n238_), .A2(KEYINPUT97), .A3(new_n246_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n239_), .A2(new_n242_), .B1(new_n236_), .B2(new_n234_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT97), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(new_n244_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n204_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n238_), .A2(KEYINPUT4), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n203_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n247_), .A2(new_n202_), .A3(new_n250_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G85gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G78gat), .B(G106gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT93), .Z(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G197gat), .A2(G204gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G197gat), .A2(G204gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT21), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT21), .ZN(new_n271_));
  AND2_X1   g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n267_), .ZN(new_n273_));
  INV_X1    g072(.A(G211gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G218gat), .ZN(new_n275_));
  INV_X1    g074(.A(G218gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT89), .B1(new_n276_), .B2(G211gat), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n270_), .A2(new_n273_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n275_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n279_), .A2(KEYINPUT21), .A3(new_n268_), .A4(new_n269_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n278_), .A2(new_n280_), .A3(KEYINPUT92), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT92), .B1(new_n278_), .B2(new_n280_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n243_), .A2(new_n245_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n266_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n278_), .A2(new_n280_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT90), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n278_), .A2(new_n280_), .A3(KEYINPUT90), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n285_), .A2(KEYINPUT29), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n266_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n265_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n287_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(new_n283_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n264_), .B(new_n295_), .C1(new_n299_), .C2(new_n266_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n300_), .A3(KEYINPUT94), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  XOR2_X1   g101(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(new_n285_), .B2(KEYINPUT29), .ZN(new_n304_));
  XOR2_X1   g103(.A(G22gat), .B(G50gat), .Z(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  INV_X1    g105(.A(new_n303_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n248_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n305_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n302_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT88), .A3(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(new_n265_), .C1(new_n288_), .C2(new_n296_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n301_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n263_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(new_n300_), .A3(new_n309_), .A4(new_n313_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G227gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(G71gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G99gat), .ZN(new_n326_));
  AND3_X1   g125(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OR3_X1    g128(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT24), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G183gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT78), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(G183gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT25), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n331_), .B(new_n336_), .C1(new_n339_), .C2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n341_), .A2(new_n348_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n329_), .A2(new_n349_), .B1(G169gat), .B2(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351_));
  OAI21_X1  g150(.A(G169gat), .B1(new_n351_), .B2(KEYINPUT79), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n332_), .A3(KEYINPUT22), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .A4(new_n333_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n354_), .A3(new_n333_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT80), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n350_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n326_), .B1(new_n347_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G15gat), .B(G43gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT81), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT30), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n347_), .A2(new_n326_), .A3(new_n359_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n360_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT83), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n366_), .A2(new_n369_), .A3(KEYINPUT82), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n244_), .B(KEYINPUT31), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n372_), .A2(new_n378_), .A3(new_n374_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT19), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G169gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n333_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n350_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n329_), .A2(new_n336_), .A3(new_n330_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n348_), .A2(KEYINPUT26), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G190gat), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n391_), .A2(new_n393_), .A3(KEYINPUT95), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT95), .B1(new_n391_), .B2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n338_), .A2(new_n342_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n389_), .B1(new_n390_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n386_), .B1(new_n398_), .B2(new_n289_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n291_), .A2(new_n347_), .A3(new_n359_), .A4(new_n292_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n385_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n347_), .A2(new_n359_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n386_), .B1(new_n293_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n395_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n340_), .A2(KEYINPUT95), .ZN(new_n412_));
  INV_X1    g211(.A(new_n396_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n390_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n414_), .A2(new_n415_), .B1(new_n350_), .B2(new_n388_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n289_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n384_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n402_), .A2(new_n408_), .A3(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n420_), .A2(KEYINPUT27), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT99), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n398_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(KEYINPUT99), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n283_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n385_), .B1(new_n425_), .B2(new_n410_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n400_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n416_), .B2(new_n417_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n384_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n407_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n410_), .A2(new_n418_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n407_), .B1(new_n431_), .B2(new_n401_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n420_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT27), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n421_), .A2(new_n430_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AND4_X1   g234(.A1(new_n262_), .A2(new_n322_), .A3(new_n382_), .A4(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n321_), .A3(new_n262_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n402_), .A2(new_n438_), .A3(new_n419_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n258_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT97), .B1(new_n248_), .B2(new_n244_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n250_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT4), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n252_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n202_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n254_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n443_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n442_), .B1(new_n452_), .B2(new_n259_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n253_), .A2(new_n254_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT33), .B1(new_n454_), .B2(new_n443_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  AOI211_X1 g255(.A(new_n456_), .B(new_n258_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n247_), .A2(new_n250_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n443_), .B1(new_n459_), .B2(new_n203_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n448_), .A2(new_n202_), .A3(new_n449_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(KEYINPUT98), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT98), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n448_), .A2(new_n464_), .A3(new_n202_), .A4(new_n449_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n433_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n453_), .B1(new_n458_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n437_), .B1(new_n467_), .B2(new_n321_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n382_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n380_), .A2(KEYINPUT84), .A3(new_n381_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n436_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT72), .B(G8gat), .ZN(new_n474_));
  INV_X1    g273(.A(G1gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT73), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n478_), .B(KEYINPUT73), .ZN(new_n483_));
  INV_X1    g282(.A(new_n481_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT71), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n491_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n487_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT76), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n498_), .B(new_n502_), .C1(KEYINPUT75), .C2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n473_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G120gat), .B(G148gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G176gat), .B(G204gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT64), .Z(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G78gat), .Z(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT67), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n533_), .A3(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT68), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT6), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT68), .B(KEYINPUT6), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(new_n540_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547_));
  INV_X1    g346(.A(G99gat), .ZN(new_n548_));
  INV_X1    g347(.A(G106gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .A4(KEYINPUT66), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n535_), .B1(new_n546_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT8), .ZN(new_n556_));
  INV_X1    g355(.A(new_n542_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n540_), .A2(new_n536_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n560_), .A2(new_n554_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n532_), .A2(new_n534_), .A3(new_n556_), .ZN(new_n562_));
  OAI22_X1  g361(.A1(new_n555_), .A2(new_n556_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT10), .B(G99gat), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n549_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT65), .B(G92gat), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(G85gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n529_), .A2(KEYINPUT9), .A3(new_n530_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n558_), .A2(new_n559_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n565_), .A2(new_n568_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n528_), .B1(new_n563_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n557_), .B1(new_n544_), .B2(new_n540_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n537_), .A2(new_n539_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(G99gat), .A3(G106gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n554_), .A3(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n532_), .A2(new_n534_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n556_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n562_), .B1(new_n554_), .B2(new_n560_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n528_), .B(new_n571_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n521_), .B1(new_n572_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT69), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT12), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n572_), .B2(new_n581_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n521_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n571_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n528_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n586_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n588_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n519_), .B1(new_n583_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n583_), .A2(new_n597_), .A3(new_n519_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n515_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n600_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(KEYINPUT13), .A3(new_n598_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n500_), .A2(new_n589_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n493_), .A2(new_n563_), .A3(new_n571_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT35), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(KEYINPUT36), .ZN(new_n619_));
  INV_X1    g418(.A(new_n614_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n606_), .A2(new_n620_), .A3(new_n607_), .A4(new_n612_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n615_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n618_), .B(KEYINPUT36), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT37), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n622_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(G231gat), .ZN(new_n633_));
  INV_X1    g432(.A(G233gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n486_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n486_), .A2(new_n635_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n528_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n590_), .A3(new_n636_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT17), .ZN(new_n643_));
  XOR2_X1   g442(.A(G127gat), .B(G155gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT16), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n642_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n643_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT74), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(KEYINPUT74), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n632_), .A2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n514_), .A2(new_n605_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n262_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n475_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n623_), .A2(new_n626_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n473_), .A2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n604_), .A2(new_n653_), .A3(new_n513_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n262_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n657_), .A2(new_n658_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n659_), .A2(new_n664_), .A3(new_n665_), .ZN(G1324gat));
  OAI21_X1  g465(.A(G8gat), .B1(new_n663_), .B2(new_n435_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT39), .ZN(new_n668_));
  INV_X1    g467(.A(new_n435_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n655_), .A2(new_n669_), .A3(new_n474_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n663_), .B2(new_n472_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT41), .Z(new_n674_));
  INV_X1    g473(.A(G15gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n472_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n655_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n655_), .A2(new_n679_), .A3(new_n321_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n663_), .B2(new_n322_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n683_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT101), .Z(G1327gat));
  INV_X1    g486(.A(new_n653_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n688_), .A2(new_n604_), .A3(new_n513_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n473_), .B2(new_n631_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n452_), .A2(new_n456_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n433_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n462_), .A2(KEYINPUT98), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n465_), .A3(new_n460_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n261_), .A2(KEYINPUT33), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n691_), .A2(new_n692_), .A3(new_n694_), .A4(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n440_), .B(new_n441_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n321_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n435_), .A2(new_n262_), .A3(new_n321_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n472_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n669_), .A2(new_n321_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n262_), .A3(new_n382_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT43), .B(new_n631_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n690_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n702_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n706_), .A2(new_n704_), .A3(new_n632_), .A4(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n689_), .B1(new_n705_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n707_), .A3(new_n632_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT102), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n708_), .A3(new_n690_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(KEYINPUT44), .A3(new_n689_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717_), .B2(new_n262_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n660_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n688_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n514_), .A2(new_n605_), .A3(new_n720_), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n721_), .A2(G29gat), .A3(new_n262_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n435_), .B(KEYINPUT105), .Z(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(KEYINPUT107), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728_));
  INV_X1    g527(.A(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n721_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT106), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n733_), .A3(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT45), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n712_), .A2(new_n737_), .A3(new_n669_), .A4(new_n716_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(G36gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n712_), .A2(new_n669_), .A3(new_n716_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT103), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT104), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  AND4_X1   g541(.A1(KEYINPUT104), .A2(new_n741_), .A3(G36gat), .A4(new_n738_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n736_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT46), .B(new_n736_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1329gat));
  NAND2_X1  g547(.A1(new_n382_), .A2(G43gat), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n721_), .A2(new_n472_), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n717_), .A2(new_n749_), .B1(G43gat), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g551(.A(G50gat), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n717_), .A2(new_n753_), .A3(new_n322_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G50gat), .B1(new_n724_), .B2(new_n321_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT108), .ZN(G1331gat));
  NOR2_X1   g556(.A1(new_n473_), .A2(new_n512_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n604_), .A3(new_n654_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT109), .Z(new_n760_));
  AOI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n656_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n605_), .A2(new_n512_), .A3(new_n653_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n661_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n262_), .A2(KEYINPUT110), .ZN(new_n765_));
  MUX2_X1   g564(.A(KEYINPUT110), .B(new_n765_), .S(G57gat), .Z(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n764_), .B2(new_n766_), .ZN(G1332gat));
  INV_X1    g566(.A(G64gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n725_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G64gat), .B1(new_n763_), .B2(new_n725_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT48), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1333gat));
  NAND3_X1  g572(.A1(new_n760_), .A2(new_n324_), .A3(new_n676_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G71gat), .B1(new_n763_), .B2(new_n472_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT49), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n760_), .A2(new_n778_), .A3(new_n321_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G78gat), .B1(new_n763_), .B2(new_n322_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT50), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n605_), .A2(new_n688_), .A3(new_n512_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n715_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n262_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n758_), .A2(new_n604_), .A3(new_n720_), .ZN(new_n787_));
  OR3_X1    g586(.A1(new_n787_), .A2(G85gat), .A3(new_n262_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT111), .Z(G1336gat));
  INV_X1    g589(.A(new_n787_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G92gat), .B1(new_n791_), .B2(new_n669_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n769_), .A2(new_n566_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n784_), .B2(new_n793_), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n785_), .B2(new_n472_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n382_), .A3(new_n564_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g597(.A(new_n549_), .B1(new_n784_), .B2(new_n321_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT52), .Z(new_n800_));
  NAND3_X1  g599(.A1(new_n791_), .A2(new_n549_), .A3(new_n321_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  INV_X1    g603(.A(G113gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n262_), .B1(new_n381_), .B2(new_n380_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n701_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n600_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n593_), .A2(new_n594_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n589_), .A2(new_n590_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n594_), .B1(new_n813_), .B2(new_n580_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n587_), .A2(KEYINPUT112), .A3(new_n595_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n521_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n812_), .A2(new_n814_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n588_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n587_), .A2(KEYINPUT55), .A3(new_n595_), .A4(new_n588_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n596_), .A2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n817_), .A2(new_n819_), .A3(new_n822_), .A4(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n519_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT114), .B(KEYINPUT56), .Z(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n825_), .B2(new_n519_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n810_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n495_), .A2(new_n496_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n501_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n510_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n508_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n833_));
  OAI22_X1  g632(.A1(new_n599_), .A2(new_n600_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n660_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n832_), .A2(new_n833_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n600_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n519_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n826_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n838_), .B(KEYINPUT58), .C1(new_n826_), .C2(new_n839_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n632_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n836_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n835_), .A2(KEYINPUT57), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n653_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n654_), .A2(new_n513_), .A3(new_n605_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT54), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n850_), .A2(KEYINPUT54), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n847_), .A2(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n809_), .B1(new_n849_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n835_), .B2(KEYINPUT57), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n837_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n519_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n519_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n587_), .A2(new_n595_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n588_), .B1(new_n861_), .B2(new_n811_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n862_), .A2(new_n816_), .B1(new_n823_), .B2(new_n596_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n820_), .B(KEYINPUT113), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n860_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n859_), .B1(new_n865_), .B2(new_n827_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n858_), .B1(new_n866_), .B2(new_n810_), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT115), .B(new_n857_), .C1(new_n867_), .C2(new_n660_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n856_), .A2(new_n868_), .A3(new_n836_), .A4(new_n844_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n653_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n852_), .A2(new_n851_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n870_), .A2(KEYINPUT116), .A3(new_n871_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n807_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n854_), .B1(new_n877_), .B2(KEYINPUT59), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n805_), .B1(new_n878_), .B2(new_n512_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n874_), .A2(KEYINPUT117), .A3(new_n875_), .A4(new_n876_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n513_), .A2(G113gat), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n804_), .B1(new_n879_), .B2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n513_), .B(new_n854_), .C1(new_n877_), .C2(KEYINPUT59), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT119), .B(new_n886_), .C1(new_n887_), .C2(new_n805_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1340gat));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n878_), .B2(new_n604_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n892_));
  AOI21_X1  g691(.A(G120gat), .B1(new_n604_), .B2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n892_), .B2(G120gat), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n881_), .A2(new_n882_), .A3(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT120), .B1(new_n891_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n881_), .A2(new_n882_), .A3(new_n894_), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n605_), .B(new_n854_), .C1(new_n877_), .C2(KEYINPUT59), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n897_), .B(new_n898_), .C1(new_n899_), .C2(new_n890_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n900_), .ZN(G1341gat));
  AND3_X1   g700(.A1(new_n878_), .A2(G127gat), .A3(new_n688_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n881_), .A2(new_n688_), .A3(new_n882_), .ZN(new_n903_));
  INV_X1    g702(.A(G127gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n903_), .A2(KEYINPUT121), .A3(new_n904_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n902_), .B1(new_n907_), .B2(new_n908_), .ZN(G1342gat));
  AND2_X1   g708(.A1(new_n878_), .A2(new_n632_), .ZN(new_n910_));
  INV_X1    g709(.A(G134gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n881_), .A2(new_n882_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n660_), .A2(new_n911_), .ZN(new_n913_));
  OAI22_X1  g712(.A1(new_n910_), .A2(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1343gat));
  NAND2_X1  g713(.A1(new_n874_), .A2(new_n875_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n676_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n769_), .A2(new_n262_), .A3(new_n322_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(new_n227_), .A3(new_n512_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G141gat), .B1(new_n918_), .B2(new_n513_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1344gat));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(G148gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n604_), .A3(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n923_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n918_), .B2(new_n605_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1345gat));
  XNOR2_X1  g726(.A(KEYINPUT61), .B(G155gat), .ZN(new_n928_));
  OR3_X1    g727(.A1(new_n918_), .A2(new_n653_), .A3(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n918_), .B2(new_n653_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n918_), .B2(new_n631_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n660_), .A2(new_n212_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n918_), .B2(new_n933_), .ZN(G1347gat));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n321_), .B1(new_n849_), .B2(new_n853_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n725_), .A2(new_n656_), .A3(new_n472_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n513_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n935_), .B1(new_n939_), .B2(new_n332_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n387_), .ZN(new_n941_));
  OAI211_X1 g740(.A(KEYINPUT62), .B(G169gat), .C1(new_n938_), .C2(new_n513_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n940_), .A2(new_n941_), .A3(new_n942_), .ZN(G1348gat));
  NOR2_X1   g742(.A1(new_n915_), .A2(new_n321_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n944_), .A2(G176gat), .A3(new_n604_), .A4(new_n937_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n333_), .B1(new_n938_), .B2(new_n605_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n945_), .A2(KEYINPUT123), .A3(new_n946_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1349gat));
  NAND2_X1  g750(.A1(new_n937_), .A2(new_n688_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n915_), .A2(new_n321_), .A3(new_n952_), .ZN(new_n953_));
  OR2_X1    g752(.A1(new_n953_), .A2(KEYINPUT124), .ZN(new_n954_));
  AOI21_X1  g753(.A(G183gat), .B1(new_n953_), .B2(KEYINPUT124), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n952_), .A2(new_n413_), .ZN(new_n956_));
  AOI22_X1  g755(.A1(new_n954_), .A2(new_n955_), .B1(new_n936_), .B2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n938_), .B2(new_n631_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n660_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n938_), .B2(new_n959_), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n725_), .A2(new_n656_), .A3(new_n322_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n916_), .A2(new_n961_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963_), .B2(new_n512_), .ZN(new_n964_));
  INV_X1    g763(.A(G197gat), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n962_), .A2(new_n965_), .A3(new_n513_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1352gat));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(G204gat), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n963_), .A2(new_n604_), .A3(new_n969_), .ZN(new_n970_));
  OAI211_X1 g769(.A(new_n968_), .B(G204gat), .C1(new_n962_), .C2(new_n605_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(G1353gat));
  AOI21_X1  g771(.A(new_n653_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n973_));
  NOR2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(KEYINPUT126), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n963_), .A2(new_n973_), .A3(new_n975_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n974_), .B(KEYINPUT126), .ZN(new_n977_));
  INV_X1    g776(.A(new_n973_), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n977_), .B1(new_n962_), .B2(new_n978_), .ZN(new_n979_));
  AND2_X1   g778(.A1(new_n976_), .A2(new_n979_), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n962_), .B2(new_n631_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n660_), .A2(new_n276_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n962_), .B2(new_n982_), .ZN(G1355gat));
endmodule


