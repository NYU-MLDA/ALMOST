//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT81), .ZN(new_n205_));
  OR3_X1    g004(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT24), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n203_), .B1(KEYINPUT80), .B2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(KEYINPUT80), .B2(new_n213_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT79), .B(G190gat), .Z(new_n217_));
  OAI211_X1 g016(.A(new_n215_), .B(new_n216_), .C1(new_n213_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n208_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT83), .B(G176gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n206_), .A2(new_n204_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n217_), .B2(G183gat), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n212_), .A2(new_n222_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT84), .B(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n230_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n234_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G1gat), .B(G29gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G85gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  OR2_X1    g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT86), .ZN(new_n256_));
  OAI22_X1  g055(.A1(new_n256_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258_));
  INV_X1    g057(.A(G141gat), .ZN(new_n259_));
  INV_X1    g058(.A(G148gat), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .A4(KEYINPUT86), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(KEYINPUT2), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(KEYINPUT2), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n257_), .B(new_n261_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT88), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n254_), .B(new_n255_), .C1(new_n266_), .C2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n259_), .A2(new_n260_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT85), .B1(new_n254_), .B2(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n254_), .A2(KEYINPUT1), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n255_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n254_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n262_), .B(new_n270_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n276_), .A2(KEYINPUT4), .A3(new_n237_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT99), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n278_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n253_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(KEYINPUT98), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(new_n237_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT4), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(KEYINPUT100), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n253_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT100), .B1(new_n281_), .B2(new_n284_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n252_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n281_), .A2(new_n284_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT100), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(new_n251_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n246_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n227_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n216_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n220_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT93), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n228_), .A2(new_n209_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n298_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G197gat), .B(G204gat), .Z(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(KEYINPUT90), .A3(KEYINPUT21), .ZN(new_n306_));
  XOR2_X1   g105(.A(G211gat), .B(G218gat), .Z(new_n307_));
  OAI22_X1  g106(.A1(new_n306_), .A2(new_n307_), .B1(KEYINPUT21), .B2(new_n305_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n306_), .A2(new_n307_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT94), .Z(new_n312_));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n313_));
  INV_X1    g112(.A(new_n310_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n230_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT20), .B1(new_n304_), .B2(new_n310_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n230_), .A2(KEYINPUT95), .A3(new_n314_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT95), .B1(new_n230_), .B2(new_n314_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n320_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n319_), .B1(new_n324_), .B2(new_n318_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G64gat), .B(G92gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT97), .ZN(new_n327_));
  XOR2_X1   g126(.A(G8gat), .B(G36gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n311_), .B(KEYINPUT94), .ZN(new_n334_));
  INV_X1    g133(.A(new_n315_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n317_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n320_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT95), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n212_), .A2(new_n222_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n227_), .A2(new_n229_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n338_), .B1(new_n341_), .B2(new_n310_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n318_), .B(new_n337_), .C1(new_n342_), .C2(new_n321_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n336_), .A2(new_n343_), .A3(new_n331_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT102), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n336_), .A2(new_n343_), .A3(KEYINPUT102), .A4(new_n331_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n333_), .A2(new_n346_), .A3(KEYINPUT27), .A4(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n336_), .A2(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n332_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n344_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n276_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G22gat), .B(G50gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n355_), .B(KEYINPUT28), .ZN(new_n360_));
  INV_X1    g159(.A(new_n358_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT92), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT92), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT89), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n314_), .B2(KEYINPUT91), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n310_), .B1(new_n276_), .B2(new_n354_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G78gat), .B(G106gat), .Z(new_n373_));
  INV_X1    g172(.A(new_n371_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n363_), .A2(new_n374_), .A3(KEYINPUT92), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n373_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n348_), .A2(new_n353_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT103), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n348_), .A2(new_n353_), .A3(KEYINPUT103), .A4(new_n378_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n296_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n279_), .A2(new_n280_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n284_), .A2(new_n385_), .A3(new_n253_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n253_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n251_), .B1(new_n283_), .B2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n293_), .A2(new_n384_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n287_), .A2(new_n288_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(KEYINPUT33), .A3(new_n251_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n389_), .A2(new_n391_), .A3(new_n344_), .A4(new_n350_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n325_), .A2(KEYINPUT32), .A3(new_n331_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n336_), .A2(new_n343_), .A3(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n294_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n378_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n378_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n399_), .A2(new_n348_), .A3(new_n353_), .A4(new_n295_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n246_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n383_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT78), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G1gat), .A2(G8gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT14), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT73), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n407_), .A3(KEYINPUT14), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G15gat), .B(G22gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G1gat), .B(G8gat), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(new_n406_), .A3(new_n408_), .A4(new_n409_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G43gat), .B(G50gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G36gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G29gat), .ZN(new_n420_));
  INV_X1    g219(.A(G29gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G36gat), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n420_), .A2(new_n422_), .A3(KEYINPUT68), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT68), .B1(new_n420_), .B2(new_n422_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n418_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n422_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT68), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n420_), .A2(new_n422_), .A3(KEYINPUT68), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n417_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT75), .B1(new_n416_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n430_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n415_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n415_), .A2(new_n433_), .A3(KEYINPUT76), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT76), .B1(new_n415_), .B2(new_n433_), .ZN(new_n437_));
  OAI22_X1  g236(.A1(new_n432_), .A2(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT77), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G229gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n437_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n415_), .A2(new_n433_), .A3(KEYINPUT76), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n416_), .A2(new_n431_), .A3(KEYINPUT75), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n434_), .B1(new_n415_), .B2(new_n433_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n439_), .A2(new_n441_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT15), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n433_), .B(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n415_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n447_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n440_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G113gat), .B(G141gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G169gat), .B(G197gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n450_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n403_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n450_), .A2(new_n455_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n458_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(KEYINPUT78), .A3(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n402_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G120gat), .B(G148gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT5), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G176gat), .B(G204gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G64gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n477_));
  XOR2_X1   g276(.A(G71gat), .B(G78gat), .Z(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n483_), .A2(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G85gat), .ZN(new_n494_));
  INV_X1    g293(.A(G92gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(KEYINPUT9), .A3(new_n486_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n489_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT64), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n489_), .A2(new_n500_), .A3(new_n493_), .A4(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n487_), .A2(new_n503_), .A3(KEYINPUT8), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n483_), .A2(new_n485_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  INV_X1    g305(.A(G99gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n491_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n504_), .B(KEYINPUT65), .C1(new_n505_), .C2(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  INV_X1    g315(.A(new_n509_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT66), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n483_), .A2(new_n485_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n508_), .A2(new_n521_), .A3(new_n509_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n487_), .A2(new_n503_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n516_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n481_), .B(new_n502_), .C1(new_n515_), .C2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G230gat), .ZN(new_n527_));
  INV_X1    g326(.A(G233gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n524_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n510_), .A2(KEYINPUT66), .B1(new_n483_), .B2(new_n485_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n533_), .B2(new_n522_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n513_), .B(new_n514_), .C1(new_n534_), .C2(new_n516_), .ZN(new_n535_));
  AOI211_X1 g334(.A(KEYINPUT12), .B(new_n481_), .C1(new_n535_), .C2(new_n502_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT12), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n502_), .B1(new_n515_), .B2(new_n525_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n481_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n531_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n539_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n530_), .B1(new_n542_), .B2(new_n526_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n474_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n544_), .A3(new_n474_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(KEYINPUT67), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n549_));
  INV_X1    g348(.A(new_n547_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(new_n551_), .A3(KEYINPUT13), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT36), .Z(new_n561_));
  OAI211_X1 g360(.A(new_n431_), .B(new_n502_), .C1(new_n515_), .C2(new_n525_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n535_), .A2(KEYINPUT69), .A3(new_n431_), .A4(new_n502_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT34), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n452_), .A2(new_n538_), .B1(new_n570_), .B2(new_n569_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n572_), .B1(new_n566_), .B2(new_n573_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n566_), .A2(new_n573_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n571_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT71), .B1(new_n580_), .B2(new_n574_), .ZN(new_n581_));
  OAI211_X1 g380(.A(KEYINPUT72), .B(new_n561_), .C1(new_n578_), .C2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n583_), .A3(new_n574_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT70), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n580_), .A2(new_n586_), .A3(new_n583_), .A4(new_n574_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n577_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n580_), .A2(KEYINPUT71), .A3(new_n574_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT72), .B1(new_n592_), .B2(new_n561_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n557_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n415_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n481_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT16), .ZN(new_n599_));
  XOR2_X1   g398(.A(G183gat), .B(G211gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n597_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  MUX2_X1   g403(.A(new_n603_), .B(KEYINPUT17), .S(new_n601_), .Z(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n597_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n580_), .A2(new_n574_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n557_), .B1(new_n607_), .B2(new_n561_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n588_), .A2(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n594_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n469_), .A2(new_n556_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G1gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n294_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n561_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT72), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n588_), .A3(new_n582_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n402_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n556_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n621_), .A2(new_n467_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n606_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n625_), .B2(new_n295_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n613_), .A2(new_n614_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n615_), .A2(new_n626_), .A3(new_n627_), .ZN(G1324gat));
  INV_X1    g427(.A(G8gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n348_), .A2(new_n353_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n611_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n630_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G8gat), .B1(new_n625_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n635_), .B(G8gat), .C1(new_n625_), .C2(new_n632_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n631_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT40), .B(new_n631_), .C1(new_n634_), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1325gat));
  INV_X1    g441(.A(new_n246_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G15gat), .B1(new_n625_), .B2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT41), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n611_), .A2(new_n240_), .A3(new_n246_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1326gat));
  OAI21_X1  g446(.A(G22gat), .B1(new_n625_), .B2(new_n378_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n611_), .A2(new_n650_), .A3(new_n399_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(G1327gat));
  NOR3_X1   g451(.A1(new_n621_), .A2(new_n606_), .A3(new_n619_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n469_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G29gat), .B1(new_n655_), .B2(new_n294_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n594_), .A2(new_n609_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n383_), .B2(new_n401_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n657_), .B(new_n661_), .C1(new_n383_), .C2(new_n401_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n606_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n622_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT44), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n295_), .A2(new_n421_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n656_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n654_), .A2(G36gat), .A3(new_n632_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n672_), .B(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n419_), .B1(new_n668_), .B2(new_n630_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n667_), .B(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G36gat), .B1(new_n679_), .B2(new_n632_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n672_), .B(new_n673_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n681_), .A3(KEYINPUT46), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n677_), .A2(new_n682_), .ZN(G1329gat));
  XNOR2_X1  g482(.A(KEYINPUT106), .B(G43gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n655_), .B2(new_n246_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n246_), .A2(G43gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n668_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1330gat));
  OR3_X1    g488(.A1(new_n654_), .A2(G50gat), .A3(new_n378_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n668_), .A2(KEYINPUT107), .A3(new_n399_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G50gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT107), .B1(new_n668_), .B2(new_n399_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(G1331gat));
  NOR2_X1   g493(.A1(new_n556_), .A2(new_n468_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n402_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(new_n610_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n294_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n620_), .A2(new_n606_), .A3(new_n695_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G57gat), .B1(new_n700_), .B2(new_n295_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n700_), .B2(new_n632_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT48), .ZN(new_n704_));
  INV_X1    g503(.A(G64gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n697_), .A2(new_n705_), .A3(new_n630_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1333gat));
  OAI21_X1  g506(.A(G71gat), .B1(new_n700_), .B2(new_n643_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT49), .ZN(new_n709_));
  INV_X1    g508(.A(G71gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n697_), .A2(new_n710_), .A3(new_n246_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1334gat));
  OAI21_X1  g511(.A(G78gat), .B1(new_n700_), .B2(new_n378_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n378_), .A2(G78gat), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT109), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n697_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n619_), .A2(new_n606_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n696_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n494_), .A3(new_n294_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n695_), .A2(new_n664_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n295_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1336gat));
  OAI21_X1  g527(.A(new_n495_), .B1(new_n721_), .B2(new_n632_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT110), .Z(new_n730_));
  NOR3_X1   g529(.A1(new_n726_), .A2(new_n495_), .A3(new_n632_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n726_), .B2(new_n643_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n246_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n733_), .B(new_n734_), .C1(new_n721_), .C2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g536(.A1(new_n722_), .A2(new_n491_), .A3(new_n399_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n378_), .B(new_n724_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n491_), .B1(new_n740_), .B2(KEYINPUT112), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT112), .B1(new_n725_), .B2(new_n399_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n739_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n724_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n663_), .A2(KEYINPUT112), .A3(new_n399_), .A4(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G106gat), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(KEYINPUT52), .A3(new_n742_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n738_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n738_), .C1(new_n744_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1339gat));
  INV_X1    g552(.A(KEYINPUT59), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n610_), .A2(new_n756_), .A3(new_n467_), .A4(new_n556_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n594_), .A2(new_n556_), .A3(new_n606_), .A4(new_n609_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT54), .B1(new_n758_), .B2(new_n468_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n619_), .A2(new_n557_), .B1(new_n588_), .B2(new_n608_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n526_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n529_), .ZN(new_n763_));
  XOR2_X1   g562(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n764_));
  NAND2_X1  g563(.A1(new_n541_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n531_), .B(KEYINPUT55), .C1(new_n536_), .C2(new_n540_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n473_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n473_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n438_), .A2(KEYINPUT77), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n448_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n440_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n453_), .A2(new_n447_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n458_), .B1(new_n774_), .B2(new_n441_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n441_), .B1(new_n439_), .B2(new_n449_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n459_), .B1(new_n454_), .B2(new_n440_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT116), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n780_), .B2(new_n462_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n547_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n761_), .B1(new_n770_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n776_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n465_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n550_), .B1(new_n785_), .B2(new_n777_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n786_), .B(KEYINPUT58), .C1(new_n768_), .C2(new_n769_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT117), .B1(new_n760_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n657_), .A2(new_n790_), .A3(new_n783_), .A4(new_n787_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n781_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n529_), .A2(new_n762_), .B1(new_n541_), .B2(new_n764_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n474_), .B1(new_n795_), .B2(new_n766_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n767_), .B2(new_n473_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT115), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n796_), .A2(KEYINPUT56), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n463_), .A2(new_n466_), .A3(new_n547_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n793_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n619_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n792_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n768_), .B1(KEYINPUT115), .B2(new_n799_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n803_), .B1(new_n808_), .B2(new_n798_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n619_), .C1(new_n809_), .C2(new_n793_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n789_), .A2(new_n791_), .A3(new_n807_), .A4(new_n810_), .ZN(new_n811_));
  AOI221_X4 g610(.A(new_n755_), .B1(new_n757_), .B2(new_n759_), .C1(new_n811_), .C2(new_n664_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n664_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n757_), .A2(new_n759_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT118), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n295_), .B(new_n643_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n754_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n807_), .B(new_n810_), .C1(new_n760_), .C2(new_n788_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n664_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n814_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n821_), .A2(new_n817_), .A3(KEYINPUT119), .A4(new_n754_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n817_), .A2(new_n754_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n819_), .A2(new_n664_), .B1(new_n759_), .B2(new_n757_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT120), .B1(new_n818_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n381_), .A2(new_n382_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n294_), .A3(new_n246_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n812_), .A2(new_n815_), .A3(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n830_), .B(new_n827_), .C1(new_n833_), .C2(new_n754_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n468_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G113gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n833_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n467_), .A2(G113gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n818_), .A2(new_n828_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n621_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n556_), .A2(KEYINPUT60), .ZN(new_n844_));
  MUX2_X1   g643(.A(KEYINPUT60), .B(new_n844_), .S(new_n840_), .Z(new_n845_));
  NAND2_X1  g644(.A1(new_n833_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(KEYINPUT121), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  INV_X1    g647(.A(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n842_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(G1341gat));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n664_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n829_), .A2(new_n834_), .A3(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n837_), .B2(new_n664_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(KEYINPUT122), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n829_), .A2(new_n657_), .A3(new_n834_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G134gat), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n619_), .A2(G134gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n837_), .B2(new_n863_), .ZN(G1343gat));
  INV_X1    g663(.A(new_n816_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n246_), .A2(new_n378_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n632_), .A2(new_n294_), .A3(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n468_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n621_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n606_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  AND3_X1   g674(.A1(new_n868_), .A2(G162gat), .A3(new_n657_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G162gat), .B1(new_n868_), .B2(new_n806_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n878_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(G1347gat));
  NAND3_X1  g680(.A1(new_n630_), .A2(new_n295_), .A3(new_n246_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n825_), .A2(new_n399_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n467_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT124), .B1(new_n884_), .B2(new_n467_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(G169gat), .A3(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n889_), .A2(new_n890_), .B1(new_n223_), .B2(new_n885_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n890_), .B2(new_n889_), .ZN(G1348gat));
  AOI21_X1  g691(.A(new_n225_), .B1(new_n883_), .B2(new_n621_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT126), .Z(new_n894_));
  NOR2_X1   g693(.A1(new_n865_), .A2(new_n399_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n882_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n896_), .A2(G176gat), .A3(new_n621_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n894_), .B1(new_n895_), .B2(new_n897_), .ZN(G1349gat));
  NOR3_X1   g697(.A1(new_n884_), .A2(new_n216_), .A3(new_n664_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n606_), .A3(new_n896_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n202_), .ZN(G1350gat));
  AOI21_X1  g700(.A(new_n203_), .B1(new_n883_), .B2(new_n657_), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT127), .Z(new_n903_));
  NAND3_X1  g702(.A1(new_n883_), .A2(new_n299_), .A3(new_n806_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  AND4_X1   g704(.A1(new_n630_), .A2(new_n816_), .A3(new_n295_), .A4(new_n866_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n468_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n621_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n606_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AND2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n911_), .B2(new_n912_), .ZN(G1354gat));
  INV_X1    g714(.A(G218gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n906_), .A2(new_n916_), .A3(new_n806_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n906_), .A2(new_n657_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1355gat));
endmodule


