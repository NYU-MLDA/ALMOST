//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT81), .B1(new_n205_), .B2(KEYINPUT25), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT83), .B1(new_n207_), .B2(KEYINPUT26), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n208_), .B(new_n211_), .C1(KEYINPUT82), .C2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT25), .B(G183gat), .Z(new_n214_));
  AOI211_X1 g013(.A(new_n206_), .B(new_n213_), .C1(KEYINPUT81), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n216_));
  INV_X1    g015(.A(new_n212_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n219_), .B(KEYINPUT23), .Z(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n220_), .B1(KEYINPUT24), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n224_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n218_), .B(new_n226_), .C1(KEYINPUT24), .C2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n223_), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT22), .B(G169gat), .Z(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  OAI221_X1 g030(.A(new_n229_), .B1(G176gat), .B2(new_n230_), .C1(new_n220_), .C2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT30), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G43gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n228_), .A2(new_n232_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT30), .ZN(new_n241_));
  OAI21_X1  g040(.A(G43gat), .B1(new_n241_), .B2(new_n237_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G99gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n239_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n204_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n239_), .A2(new_n242_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n243_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n204_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n239_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n254_), .ZN(new_n256_));
  MUX2_X1   g055(.A(new_n255_), .B(new_n256_), .S(KEYINPUT84), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT85), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n247_), .A2(new_n252_), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n258_), .B(KEYINPUT85), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G22gat), .B(G50gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT86), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT87), .ZN(new_n269_));
  OR2_X1    g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT88), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(G155gat), .B2(G162gat), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(G155gat), .A3(G162gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT89), .Z(new_n276_));
  OAI211_X1 g075(.A(new_n267_), .B(new_n269_), .C1(new_n274_), .C2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n271_), .B1(G155gat), .B2(G162gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n267_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n266_), .A2(new_n279_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT91), .B1(KEYINPUT90), .B2(KEYINPUT3), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n268_), .B2(new_n282_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n280_), .B(new_n283_), .C1(new_n268_), .C2(new_n282_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n278_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n277_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n265_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n289_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT93), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(new_n264_), .A3(new_n290_), .ZN(new_n296_));
  INV_X1    g095(.A(G228gat), .ZN(new_n297_));
  INV_X1    g096(.A(G233gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT92), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT92), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n297_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G106gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n293_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309_));
  INV_X1    g108(.A(G204gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(G197gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT94), .B(G204gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n313_), .B2(G197gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n309_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(KEYINPUT21), .C1(new_n315_), .C2(new_n314_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT96), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  OAI211_X1 g118(.A(KEYINPUT21), .B(new_n319_), .C1(new_n312_), .C2(G197gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n314_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n320_), .B(new_n309_), .C1(new_n321_), .C2(KEYINPUT21), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n287_), .A2(new_n289_), .ZN(new_n324_));
  OAI21_X1  g123(.A(G78gat), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n322_), .ZN(new_n326_));
  INV_X1    g125(.A(G78gat), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n326_), .B(new_n327_), .C1(new_n289_), .C2(new_n287_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n308_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n308_), .A3(new_n328_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n306_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  OAI22_X1  g132(.A1(new_n333_), .A2(new_n329_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n326_), .B2(new_n240_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n220_), .B1(new_n338_), .B2(new_n224_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n225_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n214_), .B(KEYINPUT98), .Z(new_n341_));
  NOR2_X1   g140(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n217_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  OAI221_X1 g143(.A(new_n339_), .B1(new_n338_), .B2(new_n340_), .C1(new_n341_), .C2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n318_), .A2(new_n322_), .A3(new_n232_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n337_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT19), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n323_), .A2(new_n233_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n345_), .A2(new_n232_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n326_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n352_), .A2(KEYINPUT20), .A3(new_n349_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT32), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G92gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT18), .B(G64gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n356_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n347_), .A2(new_n349_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n352_), .A2(KEYINPUT20), .A3(new_n354_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n349_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n287_), .A2(new_n257_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT100), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n287_), .A2(new_n255_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n374_), .B(KEYINPUT4), .C1(new_n257_), .C2(new_n287_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n369_), .A2(KEYINPUT100), .A3(new_n370_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n373_), .A2(new_n375_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n369_), .B1(new_n255_), .B2(new_n287_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n379_), .A2(new_n381_), .A3(new_n387_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n366_), .A2(new_n368_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n335_), .B1(new_n363_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n351_), .A2(new_n355_), .A3(new_n362_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n362_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT102), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n380_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n380_), .A2(new_n397_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n377_), .A3(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n388_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n390_), .A2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n390_), .A2(new_n403_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n396_), .A2(new_n402_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n263_), .B1(new_n392_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n366_), .A2(new_n362_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n395_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT27), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n389_), .A2(new_n390_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n335_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n412_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(new_n335_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n261_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n245_), .A2(new_n246_), .A3(new_n204_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n250_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n247_), .A2(new_n252_), .A3(new_n259_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(new_n413_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n407_), .A2(new_n416_), .B1(new_n418_), .B2(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  AND2_X1   g229(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n431_));
  NOR2_X1   g230(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI22_X1  g232(.A1(KEYINPUT69), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n429_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G85gat), .B(G92gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT70), .B1(new_n437_), .B2(KEYINPUT8), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT8), .ZN(new_n440_));
  AOI211_X1 g239(.A(new_n439_), .B(new_n440_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n429_), .A2(KEYINPUT68), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n433_), .A2(new_n434_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n442_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n438_), .A2(new_n441_), .A3(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT10), .B(G99gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT65), .ZN(new_n451_));
  INV_X1    g250(.A(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT9), .ZN(new_n454_));
  INV_X1    g253(.A(G85gat), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  NAND3_X1  g257(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n457_), .A2(KEYINPUT66), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n458_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n460_), .B(new_n463_), .C1(KEYINPUT66), .C2(new_n457_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n453_), .A2(new_n464_), .A3(new_n446_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n449_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G29gat), .B(G36gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G43gat), .B(G50gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n469_), .B(KEYINPUT15), .Z(new_n470_));
  OR2_X1    g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G232gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT34), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n466_), .A2(new_n469_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n472_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n471_), .A2(new_n476_), .B1(KEYINPUT73), .B2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(KEYINPUT73), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  XOR2_X1   g280(.A(G190gat), .B(G218gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(G134gat), .B(G162gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n479_), .B(new_n480_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n485_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT37), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n493_), .A3(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT74), .B(G22gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G15gat), .ZN(new_n497_));
  INV_X1    g296(.A(G1gat), .ZN(new_n498_));
  INV_X1    g297(.A(G8gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G1gat), .B(G8gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G57gat), .ZN(new_n504_));
  INV_X1    g303(.A(G64gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G57gat), .A2(G64gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT11), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G71gat), .B(G78gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT11), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(new_n512_), .A3(new_n507_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n503_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G231gat), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n298_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n298_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G183gat), .B(G211gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G127gat), .B(G155gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n519_), .B(new_n520_), .C1(KEYINPUT17), .C2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(KEYINPUT71), .A3(KEYINPUT17), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT76), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n426_), .A2(new_n495_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n437_), .A2(KEYINPUT8), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n439_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n448_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n437_), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n453_), .A2(new_n446_), .A3(new_n464_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n516_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n516_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n516_), .A2(KEYINPUT71), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n514_), .A2(new_n543_), .A3(new_n515_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n542_), .A2(KEYINPUT12), .A3(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n449_), .B2(new_n465_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n538_), .C1(new_n540_), .C2(KEYINPUT12), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G230gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT64), .ZN(new_n549_));
  MUX2_X1   g348(.A(new_n541_), .B(new_n547_), .S(new_n549_), .Z(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT72), .B(G204gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT5), .B(G176gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n556_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(KEYINPUT13), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n502_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n501_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n469_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n503_), .A2(new_n469_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(KEYINPUT77), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n503_), .A2(KEYINPUT77), .A3(new_n469_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n503_), .A2(new_n470_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n565_), .A2(new_n566_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n571_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT78), .ZN(new_n579_));
  XOR2_X1   g378(.A(G169gat), .B(G197gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(G141gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT79), .B(G113gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n579_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n573_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT80), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n563_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n531_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n498_), .A3(new_n413_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT103), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n426_), .A2(new_n491_), .A3(new_n530_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n590_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n498_), .B1(new_n597_), .B2(new_n413_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n592_), .A2(KEYINPUT103), .A3(new_n593_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n599_), .B(new_n600_), .C1(new_n593_), .C2(new_n592_), .ZN(G1324gat));
  INV_X1    g400(.A(new_n417_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G8gat), .B1(new_n596_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n591_), .A2(new_n499_), .A3(new_n417_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n605_), .A2(KEYINPUT40), .A3(new_n606_), .A4(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1325gat));
  OAI21_X1  g413(.A(G15gat), .B1(new_n596_), .B2(new_n424_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT41), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n591_), .A2(new_n203_), .A3(new_n263_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n591_), .A2(new_n619_), .A3(new_n335_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n332_), .A2(new_n334_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G22gat), .B1(new_n596_), .B2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(KEYINPUT42), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(KEYINPUT42), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT105), .ZN(G1327gat));
  INV_X1    g425(.A(new_n491_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n426_), .A2(new_n627_), .A3(new_n529_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n590_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n413_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n391_), .A2(new_n363_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n409_), .A2(new_n405_), .A3(new_n393_), .A4(new_n404_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n402_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n632_), .B(new_n621_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n416_), .A2(new_n424_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n425_), .A2(new_n418_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT43), .B1(new_n638_), .B2(new_n495_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  INV_X1    g439(.A(new_n495_), .ZN(new_n641_));
  AOI211_X1 g440(.A(new_n640_), .B(new_n641_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(KEYINPUT44), .A3(new_n590_), .A4(new_n530_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n426_), .B2(new_n641_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(KEYINPUT43), .A3(new_n495_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n590_), .A3(new_n646_), .A4(new_n530_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n644_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n413_), .A2(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n631_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n649_), .A3(new_n417_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT106), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n644_), .A2(new_n649_), .A3(new_n655_), .A4(new_n417_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(G36gat), .A3(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n629_), .A2(G36gat), .A3(new_n602_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT45), .Z(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n659_), .A3(KEYINPUT46), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  NAND3_X1  g463(.A1(new_n650_), .A2(G43gat), .A3(new_n263_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n236_), .B1(new_n629_), .B2(new_n424_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT107), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g468(.A(G50gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n630_), .A2(new_n670_), .A3(new_n335_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n650_), .A2(new_n335_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n670_), .ZN(G1331gat));
  INV_X1    g472(.A(new_n563_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n589_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n531_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G57gat), .B1(new_n677_), .B2(new_n413_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n595_), .A2(new_n676_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n679_), .A2(new_n504_), .A3(new_n414_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1332gat));
  NAND3_X1  g480(.A1(new_n677_), .A2(new_n505_), .A3(new_n417_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n595_), .A2(new_n417_), .A3(new_n676_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(G64gat), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G64gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g487(.A(G71gat), .B1(new_n679_), .B2(new_n424_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT49), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n424_), .A2(G71gat), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT110), .Z(new_n692_));
  NAND2_X1  g491(.A1(new_n677_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1334gat));
  NAND3_X1  g493(.A1(new_n677_), .A2(new_n327_), .A3(new_n335_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G78gat), .B1(new_n679_), .B2(new_n621_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT111), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT111), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT50), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT50), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n695_), .B1(new_n700_), .B2(new_n701_), .ZN(G1335gat));
  NAND2_X1  g501(.A1(new_n628_), .A2(new_n676_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n455_), .B1(new_n703_), .B2(new_n414_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n645_), .A2(new_n530_), .A3(new_n646_), .A4(new_n676_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n413_), .A2(G85gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(new_n456_), .B1(new_n703_), .B2(new_n602_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n417_), .A2(G92gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n705_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(G1337gat));
  OAI21_X1  g511(.A(G99gat), .B1(new_n705_), .B2(new_n424_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n263_), .A2(new_n451_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n703_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g515(.A(KEYINPUT52), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n705_), .A2(new_n621_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G106gat), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n717_), .B(G106gat), .C1(new_n705_), .C2(new_n621_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n335_), .A2(new_n452_), .ZN(new_n722_));
  OAI22_X1  g521(.A1(new_n719_), .A2(new_n721_), .B1(new_n703_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g523(.A(KEYINPUT54), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n492_), .A2(new_n589_), .A3(new_n494_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n563_), .A2(new_n530_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NOR4_X1   g528(.A1(new_n726_), .A2(KEYINPUT54), .A3(new_n563_), .A4(new_n530_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n558_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  INV_X1    g532(.A(new_n549_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n547_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT112), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n547_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n547_), .A2(new_n734_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n739_), .B(new_n733_), .C1(new_n547_), .C2(new_n734_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .A4(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(KEYINPUT56), .A3(new_n555_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n743_), .A3(new_n555_), .ZN(new_n744_));
  OR2_X1    g543(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n743_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n741_), .A2(new_n743_), .A3(new_n555_), .A4(new_n745_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n732_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT80), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n587_), .B(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n576_), .A2(new_n572_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n583_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n559_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n627_), .B1(new_n749_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT115), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT57), .ZN(new_n760_));
  INV_X1    g559(.A(new_n742_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n555_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n558_), .B(new_n756_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n742_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(KEYINPUT58), .A3(new_n558_), .A4(new_n756_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n768_), .A3(new_n495_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n758_), .A2(KEYINPUT115), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n760_), .A2(new_n769_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n731_), .B1(new_n772_), .B2(new_n530_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n418_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n424_), .A2(new_n414_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n773_), .A2(new_n774_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G113gat), .B1(new_n777_), .B2(new_n675_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n731_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n758_), .A2(KEYINPUT115), .A3(new_n770_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n758_), .B2(KEYINPUT115), .ZN(new_n781_));
  INV_X1    g580(.A(new_n769_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n783_), .B2(new_n529_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT59), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(new_n418_), .A3(new_n775_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n773_), .B2(KEYINPUT116), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n777_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n589_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n778_), .B1(new_n792_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  INV_X1    g593(.A(G120gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n791_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n563_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n674_), .B2(KEYINPUT60), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT117), .B1(new_n795_), .B2(KEYINPUT60), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n777_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n798_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n794_), .B1(new_n797_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n674_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n806_));
  OAI221_X1 g605(.A(KEYINPUT118), .B1(new_n801_), .B2(new_n803_), .C1(new_n806_), .C2(new_n795_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1341gat));
  AOI21_X1  g607(.A(G127gat), .B1(new_n777_), .B2(new_n529_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n530_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g610(.A(G134gat), .B1(new_n777_), .B2(new_n491_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT119), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT120), .B(G134gat), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n641_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n796_), .B2(new_n815_), .ZN(G1343gat));
  NOR2_X1   g615(.A1(new_n263_), .A2(new_n621_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n784_), .A2(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n818_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n675_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n563_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT121), .B(G148gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1345gat));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n529_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT61), .B(G155gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1346gat));
  AOI21_X1  g626(.A(G162gat), .B1(new_n819_), .B2(new_n491_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n495_), .A2(G162gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n819_), .B2(new_n829_), .ZN(G1347gat));
  NOR2_X1   g629(.A1(new_n773_), .A2(new_n335_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n602_), .A2(new_n413_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n424_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n675_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT122), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n221_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT62), .Z(new_n838_));
  AND3_X1   g637(.A1(new_n831_), .A2(KEYINPUT123), .A3(new_n834_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT123), .B1(new_n831_), .B2(new_n834_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n589_), .A2(new_n230_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n838_), .B1(new_n841_), .B2(new_n842_), .ZN(G1348gat));
  NAND2_X1  g642(.A1(new_n831_), .A2(new_n834_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n844_), .A2(new_n222_), .A3(new_n674_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n831_), .A2(KEYINPUT123), .A3(new_n834_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n674_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT124), .B1(new_n849_), .B2(G176gat), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n851_), .B(new_n222_), .C1(new_n841_), .C2(new_n674_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n845_), .B1(new_n850_), .B2(new_n852_), .ZN(G1349gat));
  NOR2_X1   g652(.A1(new_n841_), .A2(new_n530_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n831_), .A2(new_n529_), .A3(new_n834_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n854_), .A2(new_n341_), .B1(new_n205_), .B2(new_n855_), .ZN(G1350gat));
  OAI21_X1  g655(.A(G190gat), .B1(new_n841_), .B2(new_n641_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n491_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n344_), .B2(new_n858_), .ZN(G1351gat));
  NAND3_X1  g658(.A1(new_n784_), .A2(new_n817_), .A3(new_n832_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n675_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g662(.A1(new_n860_), .A2(new_n674_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n313_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n310_), .B2(new_n864_), .ZN(G1353gat));
  NAND2_X1  g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n861_), .A2(new_n529_), .A3(new_n867_), .A4(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n860_), .B2(new_n530_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT125), .B(KEYINPUT126), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1354gat));
  AOI21_X1  g673(.A(KEYINPUT127), .B1(new_n861_), .B2(new_n491_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT127), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n860_), .A2(new_n876_), .A3(new_n627_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(G218gat), .A3(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n495_), .A2(G218gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n861_), .B2(new_n879_), .ZN(G1355gat));
endmodule


