//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT8), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT68), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT67), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n217_), .A2(new_n213_), .A3(new_n214_), .A4(KEYINPUT67), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n211_), .A2(new_n212_), .A3(new_n216_), .A4(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n204_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n209_), .A3(new_n218_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n224_), .A2(new_n204_), .A3(new_n222_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G85gat), .ZN(new_n229_));
  INV_X1    g028(.A(G92gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT9), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n221_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n232_), .A2(new_n209_), .A3(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n236_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n214_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n228_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n235_), .A2(new_n237_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT64), .ZN(new_n244_));
  AOI21_X1  g043(.A(G106gat), .B1(new_n244_), .B2(new_n238_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n232_), .A2(new_n209_), .A3(new_n233_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT66), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n227_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n245_), .B2(new_n246_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n234_), .A2(new_n241_), .A3(new_n228_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT69), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n226_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G29gat), .B(G36gat), .Z(new_n253_));
  XOR2_X1   g052(.A(G43gat), .B(G50gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT15), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n203_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n223_), .A2(new_n225_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT69), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT69), .B1(new_n249_), .B2(new_n250_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(KEYINPUT76), .A3(new_n256_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n250_), .B(new_n249_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n255_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G232gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT75), .B(KEYINPUT35), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n258_), .A2(new_n263_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n271_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n252_), .A2(new_n257_), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n275_), .B(KEYINPUT78), .Z(new_n279_));
  INV_X1    g078(.A(new_n272_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n279_), .B(new_n280_), .C1(new_n265_), .C2(new_n264_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(KEYINPUT77), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G134gat), .B(G162gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT36), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n282_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT77), .A3(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(KEYINPUT36), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n277_), .B2(new_n283_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n202_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  AOI211_X1 g096(.A(KEYINPUT37), .B(new_n295_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G127gat), .B(G155gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT16), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G183gat), .B(G211gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT17), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT81), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G64gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n310_));
  XOR2_X1   g109(.A(G71gat), .B(G78gat), .Z(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n308_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT79), .B(G8gat), .ZN(new_n317_));
  INV_X1    g116(.A(G1gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT14), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT80), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G15gat), .B(G22gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G8gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n320_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n316_), .A2(new_n327_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n316_), .A2(new_n327_), .B1(new_n305_), .B2(new_n304_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n299_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n332_));
  OR2_X1    g131(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n264_), .A2(new_n315_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT70), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n335_), .C1(new_n264_), .C2(new_n315_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n315_), .A2(KEYINPUT12), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n264_), .A2(new_n315_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n262_), .A2(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n315_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n259_), .A2(new_n347_), .A3(new_n250_), .A4(new_n249_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n336_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G120gat), .B(G148gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(G176gat), .B(G204gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n346_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT72), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT72), .B1(new_n358_), .B2(new_n359_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n332_), .B(new_n333_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n364_), .A2(KEYINPUT73), .A3(KEYINPUT13), .A4(new_n360_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n331_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n327_), .A2(new_n255_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G229gat), .A2(G233gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n325_), .A2(new_n256_), .A3(new_n326_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G113gat), .B(G141gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT82), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n375_), .B(KEYINPUT83), .Z(new_n376_));
  XNOR2_X1  g175(.A(G169gat), .B(G197gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n325_), .A2(new_n326_), .A3(new_n265_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n370_), .B1(new_n369_), .B2(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n373_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n369_), .A2(new_n380_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n370_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n378_), .B1(new_n385_), .B2(new_n372_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n368_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n379_), .B1(new_n373_), .B2(new_n381_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n372_), .A3(new_n378_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT84), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G127gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(G134gat), .ZN(new_n393_));
  INV_X1    g192(.A(G134gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(G127gat), .ZN(new_n395_));
  INV_X1    g194(.A(G113gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(G120gat), .ZN(new_n397_));
  INV_X1    g196(.A(G120gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(G113gat), .ZN(new_n399_));
  OAI22_X1  g198(.A1(new_n393_), .A2(new_n395_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G127gat), .B(G134gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n403_), .A3(KEYINPUT88), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(KEYINPUT31), .Z(new_n408_));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G169gat), .A2(G176gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT22), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G169gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(G176gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G169gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT22), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n417_), .B2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n414_), .B(new_n415_), .C1(new_n421_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT24), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(new_n422_), .A3(new_n420_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n427_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT25), .B(G183gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n415_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(new_n431_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n425_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT30), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(G15gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G71gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G99gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n437_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT86), .B(G43gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n408_), .B1(new_n447_), .B2(KEYINPUT89), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT87), .B1(new_n408_), .B2(KEYINPUT89), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT3), .ZN(new_n454_));
  NOR4_X1   g253(.A1(new_n454_), .A2(KEYINPUT92), .A3(G141gat), .A4(G148gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(G141gat), .A2(G148gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT3), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT93), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT2), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n460_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n463_));
  OAI22_X1  g262(.A1(new_n455_), .A2(new_n458_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n453_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G141gat), .ZN(new_n469_));
  INV_X1    g268(.A(G148gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n457_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n454_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT3), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n459_), .A2(new_n461_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT93), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n465_), .B(KEYINPUT94), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n474_), .A2(new_n478_), .A3(new_n479_), .A4(KEYINPUT95), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G155gat), .A2(G162gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n468_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n456_), .B1(KEYINPUT90), .B2(new_n459_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(KEYINPUT90), .B2(new_n456_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n488_));
  OR3_X1    g287(.A1(new_n481_), .A2(new_n488_), .A3(KEYINPUT1), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n483_), .B1(KEYINPUT1), .B2(new_n481_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n481_), .B2(KEYINPUT1), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n400_), .A2(new_n403_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n485_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n485_), .A2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n407_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT101), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT101), .ZN(new_n500_));
  AOI211_X1 g299(.A(new_n500_), .B(new_n407_), .C1(new_n485_), .C2(new_n493_), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT4), .B(new_n496_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n493_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n484_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n474_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n453_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n504_), .B1(new_n507_), .B2(new_n480_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(new_n407_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n503_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n502_), .A2(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n503_), .B(new_n496_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT102), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n500_), .B1(new_n508_), .B2(new_n407_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n497_), .A2(KEYINPUT101), .A3(new_n498_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n495_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT102), .B1(new_n518_), .B2(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n512_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G29gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G85gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT0), .B(G57gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G8gat), .B(G36gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT18), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G64gat), .B(G92gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n532_));
  NOR2_X1   g331(.A1(G197gat), .A2(G204gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT96), .B(G197gat), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(G204gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G211gat), .B(G218gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT21), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(KEYINPUT96), .A2(G197gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(KEYINPUT96), .A2(G197gat), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n541_), .A2(new_n542_), .A3(G204gat), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n537_), .B1(G197gat), .B2(G204gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n536_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(G204gat), .B1(new_n541_), .B2(new_n542_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n533_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT21), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n539_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n532_), .B1(new_n550_), .B2(new_n436_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G226gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(G204gat), .ZN(new_n556_));
  OR2_X1    g355(.A1(KEYINPUT96), .A2(G197gat), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n540_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n537_), .B1(new_n558_), .B2(new_n533_), .ZN(new_n559_));
  INV_X1    g358(.A(G218gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G211gat), .ZN(new_n561_));
  INV_X1    g360(.A(G211gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(G218gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n557_), .A2(new_n556_), .A3(new_n540_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n565_), .B2(new_n544_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n559_), .A2(new_n566_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n414_), .A2(new_n415_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G169gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n420_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n429_), .A2(new_n430_), .B1(new_n433_), .B2(new_n415_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n427_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT98), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT98), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n427_), .A2(new_n411_), .A3(new_n575_), .A4(new_n413_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(new_n571_), .A3(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n551_), .A2(new_n555_), .A3(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n420_), .B(new_n419_), .C1(new_n569_), .C2(new_n418_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n568_), .A2(new_n580_), .B1(new_n572_), .B2(new_n428_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n532_), .B1(new_n581_), .B2(new_n567_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n571_), .A2(new_n577_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n550_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n555_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n531_), .B1(new_n579_), .B2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n567_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT20), .B1(new_n550_), .B2(new_n436_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n554_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n551_), .A2(new_n555_), .A3(new_n578_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n530_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(KEYINPUT99), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT27), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n589_), .A2(new_n594_), .A3(new_n530_), .A4(new_n590_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n555_), .B1(new_n551_), .B2(new_n578_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n587_), .A2(new_n588_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n555_), .B2(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT27), .B(new_n591_), .C1(new_n599_), .C2(new_n530_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G228gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(G78gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n214_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G22gat), .B(G50gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT28), .B1(new_n497_), .B2(KEYINPUT29), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT28), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n508_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n550_), .B1(new_n508_), .B2(new_n610_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n613_), .A3(new_n611_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n607_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n607_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n513_), .A2(new_n514_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n518_), .A2(KEYINPUT102), .A3(new_n503_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n512_), .A3(new_n524_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n526_), .A2(new_n601_), .A3(new_n620_), .A4(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT103), .ZN(new_n626_));
  INV_X1    g425(.A(new_n619_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n617_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n596_), .A2(new_n600_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n624_), .A4(new_n526_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n624_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n592_), .A2(new_n595_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n592_), .A2(KEYINPUT100), .A3(new_n595_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n524_), .A2(KEYINPUT33), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n502_), .B2(new_n511_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n503_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n502_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n524_), .B1(new_n518_), .B2(new_n643_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n623_), .A2(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n635_), .A2(new_n640_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n589_), .A2(new_n590_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n530_), .A2(KEYINPUT32), .ZN(new_n650_));
  MUX2_X1   g449(.A(new_n599_), .B(new_n649_), .S(new_n650_), .Z(new_n651_));
  AND3_X1   g450(.A1(new_n623_), .A2(new_n512_), .A3(new_n524_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n524_), .B1(new_n623_), .B2(new_n512_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n620_), .B1(new_n648_), .B2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n452_), .B1(new_n633_), .B2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n620_), .A2(new_n629_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n652_), .A2(new_n653_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n451_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n391_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n367_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n658_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n318_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n656_), .A2(new_n659_), .ZN(new_n666_));
  AND4_X1   g465(.A1(KEYINPUT77), .A2(new_n277_), .A3(new_n283_), .A4(new_n288_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n288_), .B1(new_n291_), .B2(KEYINPUT77), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n296_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n293_), .A2(KEYINPUT104), .A3(new_n296_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n666_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n330_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n366_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n391_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n674_), .A2(new_n675_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n318_), .B1(new_n679_), .B2(new_n662_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n665_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n664_), .B2(new_n663_), .ZN(G1324gat));
  INV_X1    g481(.A(G8gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n679_), .B2(new_n629_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT39), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n661_), .A2(new_n629_), .A3(new_n317_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g487(.A(new_n439_), .B1(new_n679_), .B2(new_n451_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT41), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n661_), .A2(new_n439_), .A3(new_n451_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1326gat));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n679_), .B2(new_n620_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n661_), .A2(new_n693_), .A3(new_n620_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1327gat));
  NOR2_X1   g497(.A1(new_n678_), .A2(new_n330_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  INV_X1    g499(.A(new_n299_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n666_), .B2(new_n701_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT43), .B(new_n299_), .C1(new_n656_), .C2(new_n659_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n699_), .B(KEYINPUT44), .C1(new_n702_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n658_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n366_), .A2(new_n673_), .A3(new_n330_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n660_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n658_), .A2(G29gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT46), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n629_), .A3(new_n707_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(KEYINPUT106), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n706_), .A2(new_n719_), .A3(new_n629_), .A4(new_n707_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n717_), .A2(KEYINPUT106), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(KEYINPUT107), .A3(G36gat), .A4(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n601_), .A2(G36gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT108), .B1(new_n711_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n710_), .A2(new_n660_), .A3(new_n729_), .A4(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(KEYINPUT45), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(KEYINPUT45), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n732_), .A2(new_n733_), .B1(new_n714_), .B2(KEYINPUT46), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n715_), .B1(new_n725_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n715_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n737_), .B(new_n734_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1329gat));
  OAI21_X1  g538(.A(G43gat), .B1(new_n708_), .B2(new_n452_), .ZN(new_n740_));
  INV_X1    g539(.A(G43gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n451_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n711_), .B2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT47), .Z(G1330gat));
  OR3_X1    g543(.A1(new_n711_), .A2(G50gat), .A3(new_n628_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n706_), .A2(new_n620_), .A3(new_n707_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT110), .B1(new_n746_), .B2(G50gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n366_), .A2(new_n391_), .ZN(new_n750_));
  OR3_X1    g549(.A1(new_n674_), .A2(new_n675_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(G57gat), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n658_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n677_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(new_n366_), .A3(new_n330_), .A4(new_n299_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n658_), .B1(new_n755_), .B2(KEYINPUT111), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(KEYINPUT111), .B2(new_n755_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n753_), .B1(new_n757_), .B2(new_n752_), .ZN(G1332gat));
  OAI21_X1  g557(.A(G64gat), .B1(new_n751_), .B2(new_n601_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT48), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n601_), .A2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n755_), .B2(new_n761_), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n751_), .B2(new_n452_), .ZN(new_n763_));
  XOR2_X1   g562(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n452_), .A2(G71gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n755_), .B2(new_n766_), .ZN(G1334gat));
  OAI21_X1  g566(.A(G78gat), .B1(new_n751_), .B2(new_n628_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT50), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n620_), .A2(new_n603_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n755_), .B2(new_n770_), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n676_), .A2(new_n330_), .A3(new_n673_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n754_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n662_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n702_), .A2(new_n703_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n775_), .A2(new_n330_), .A3(new_n750_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n662_), .A2(new_n229_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n774_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT114), .ZN(G1336gat));
  NAND3_X1  g580(.A1(new_n773_), .A2(new_n230_), .A3(new_n629_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n778_), .A2(new_n629_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n230_), .ZN(G1337gat));
  AOI21_X1  g583(.A(new_n213_), .B1(new_n778_), .B2(new_n451_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n773_), .B(new_n451_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OR3_X1    g587(.A1(new_n785_), .A2(KEYINPUT51), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n785_), .B2(new_n788_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1338gat));
  NAND3_X1  g590(.A1(new_n773_), .A2(new_n214_), .A3(new_n620_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n776_), .A2(new_n620_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G106gat), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT52), .B(new_n214_), .C1(new_n776_), .C2(new_n620_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g597(.A1(new_n451_), .A2(new_n662_), .A3(new_n657_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n367_), .A2(new_n391_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT54), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n367_), .A2(new_n803_), .A3(new_n391_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n338_), .B1(new_n348_), .B2(new_n335_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n339_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n345_), .B(KEYINPUT55), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n812_));
  NAND2_X1  g611(.A1(new_n346_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n340_), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n345_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n345_), .A2(new_n348_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n336_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n811_), .A2(new_n813_), .A3(new_n814_), .A4(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n357_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT119), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n817_), .A2(new_n820_), .A3(KEYINPUT56), .A4(new_n357_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n817_), .A2(new_n357_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI211_X1 g625(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n817_), .C2(new_n357_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n822_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n369_), .A2(new_n384_), .A3(new_n371_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n378_), .B1(new_n383_), .B2(new_n370_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n382_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n359_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n806_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n824_), .A2(new_n825_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT120), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n824_), .A2(new_n823_), .A3(new_n825_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n819_), .A4(new_n821_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n832_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n833_), .A2(new_n701_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n831_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n387_), .A2(new_n390_), .A3(new_n359_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT118), .B1(new_n817_), .B2(new_n357_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(KEYINPUT56), .ZN(new_n844_));
  AOI211_X1 g643(.A(KEYINPUT118), .B(new_n825_), .C1(new_n817_), .C2(new_n357_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n671_), .A2(new_n672_), .A3(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n847_), .A2(new_n848_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n846_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n330_), .B1(new_n840_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n805_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI211_X1 g656(.A(KEYINPUT123), .B(new_n330_), .C1(new_n840_), .C2(new_n854_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n800_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n802_), .A2(new_n804_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n853_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n846_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n839_), .A2(new_n701_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT58), .B1(new_n837_), .B2(new_n838_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n863_), .B(new_n864_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n330_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n840_), .A2(new_n854_), .A3(KEYINPUT122), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n862_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT59), .B1(new_n871_), .B2(new_n799_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT124), .B(new_n800_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n391_), .A2(new_n396_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n861_), .A2(new_n872_), .A3(new_n873_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n869_), .A2(new_n870_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n805_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n799_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n396_), .B1(new_n879_), .B2(new_n391_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT125), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n875_), .A2(new_n880_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1340gat));
  INV_X1    g684(.A(new_n879_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n398_), .B1(new_n676_), .B2(KEYINPUT60), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n886_), .B(new_n887_), .C1(KEYINPUT60), .C2(new_n398_), .ZN(new_n888_));
  AND4_X1   g687(.A1(new_n366_), .A2(new_n861_), .A3(new_n872_), .A4(new_n873_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n398_), .ZN(G1341gat));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n392_), .A3(new_n330_), .ZN(new_n891_));
  AND4_X1   g690(.A1(new_n330_), .A2(new_n861_), .A3(new_n872_), .A4(new_n873_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n392_), .ZN(G1342gat));
  OR3_X1    g692(.A1(new_n879_), .A2(G134gat), .A3(new_n673_), .ZN(new_n894_));
  AND4_X1   g693(.A1(new_n701_), .A2(new_n861_), .A3(new_n872_), .A4(new_n873_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n394_), .ZN(G1343gat));
  NAND4_X1  g695(.A1(new_n877_), .A2(new_n662_), .A3(new_n452_), .A4(new_n630_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n391_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n469_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n676_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT126), .B(G148gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n897_), .A2(new_n675_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  OAI21_X1  g704(.A(G162gat), .B1(new_n897_), .B2(new_n299_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n673_), .A2(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n897_), .B2(new_n907_), .ZN(G1347gat));
  NOR4_X1   g707(.A1(new_n452_), .A2(new_n662_), .A3(new_n620_), .A4(new_n601_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910_), .B2(new_n391_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n912_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n910_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n569_), .A3(new_n677_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n913_), .A2(new_n914_), .A3(new_n916_), .ZN(G1348gat));
  AOI21_X1  g716(.A(G176gat), .B1(new_n915_), .B2(new_n366_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n877_), .A2(new_n909_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n676_), .A2(new_n420_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1349gat));
  AOI21_X1  g720(.A(G183gat), .B1(new_n919_), .B2(new_n330_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n675_), .A2(new_n429_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n915_), .B2(new_n923_), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n910_), .B2(new_n299_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n430_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n673_), .A2(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n925_), .B1(new_n910_), .B2(new_n927_), .ZN(G1351gat));
  NAND3_X1  g727(.A1(new_n452_), .A2(new_n620_), .A3(new_n629_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n871_), .A2(new_n662_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n677_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n366_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g733(.A(new_n675_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n930_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT127), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n936_), .B(new_n938_), .Z(G1354gat));
  NOR2_X1   g738(.A1(new_n673_), .A2(G218gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n930_), .A2(new_n940_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n930_), .A2(new_n701_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n560_), .ZN(G1355gat));
endmodule


