//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n844_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT12), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  OAI22_X1  g009(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(KEYINPUT66), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT8), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT66), .B1(new_n212_), .B2(new_n213_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n213_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n226_), .A2(new_n227_), .A3(KEYINPUT9), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(G92gat), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n209_), .A2(new_n210_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n224_), .A2(new_n225_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n221_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n217_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G78gat), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n203_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n221_), .B(new_n232_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n241_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n202_), .A2(KEYINPUT12), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n246_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n243_), .A2(new_n244_), .A3(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n242_), .A2(new_n247_), .A3(new_n248_), .A4(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n218_), .A2(new_n219_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT8), .A3(new_n214_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n254_), .A2(new_n241_), .A3(new_n221_), .A4(new_n232_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n245_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n248_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n243_), .A2(KEYINPUT67), .A3(new_n244_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G120gat), .B(G148gat), .ZN(new_n260_));
  INV_X1    g059(.A(G204gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT5), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n251_), .A2(new_n259_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT70), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n251_), .A2(new_n259_), .A3(new_n268_), .A4(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n265_), .B(KEYINPUT69), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n251_), .A2(new_n259_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n270_), .A2(new_n271_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n271_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT13), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G29gat), .B(G36gat), .ZN(new_n281_));
  INV_X1    g080(.A(G43gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G50gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(G43gat), .ZN(new_n285_));
  INV_X1    g084(.A(G50gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289_));
  INV_X1    g088(.A(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT14), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G8gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(KEYINPUT79), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n284_), .A2(new_n287_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n295_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n295_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G229gat), .A2(G233gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n284_), .A2(new_n287_), .A3(KEYINPUT15), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT15), .B1(new_n284_), .B2(new_n287_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n295_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n304_), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G113gat), .B(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G169gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G197gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n306_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n306_), .B2(new_n310_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n280_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G113gat), .ZN(new_n323_));
  INV_X1    g122(.A(G120gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT30), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n327_), .A2(new_n329_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n312_), .A2(new_n264_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT23), .ZN(new_n334_));
  INV_X1    g133(.A(G183gat), .ZN(new_n335_));
  INV_X1    g134(.A(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n332_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G169gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(G176gat), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n334_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT81), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n332_), .A2(new_n343_), .A3(new_n342_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT80), .ZN(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT26), .B(G190gat), .Z(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(KEYINPUT25), .B2(new_n335_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n347_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n341_), .B1(new_n346_), .B2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G15gat), .B(G43gat), .Z(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT31), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n355_), .B(new_n357_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n330_), .A2(new_n331_), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT82), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT83), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n364_), .B(new_n365_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n367_), .A2(new_n370_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n363_), .B(KEYINPUT3), .Z(new_n373_));
  XOR2_X1   g172(.A(new_n365_), .B(KEYINPUT2), .Z(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT29), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT88), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT21), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT87), .B1(new_n314_), .B2(G204gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(new_n261_), .A3(G197gat), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n382_), .A2(new_n384_), .B1(new_n314_), .B2(G204gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n380_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n314_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n261_), .A2(G197gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT85), .B1(new_n314_), .B2(G204gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT21), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT86), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n386_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n385_), .A2(new_n381_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n380_), .A2(new_n395_), .A3(KEYINPUT89), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n380_), .A2(new_n395_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n377_), .A2(new_n378_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n378_), .B1(new_n377_), .B2(new_n400_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OR3_X1    g203(.A1(new_n401_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n376_), .A2(KEYINPUT29), .A3(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n376_), .B2(KEYINPUT29), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G22gat), .B(G50gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n411_), .A3(new_n409_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n405_), .B(new_n406_), .C1(new_n416_), .C2(KEYINPUT90), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n405_), .A2(new_n406_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(KEYINPUT90), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n376_), .A2(new_n431_), .A3(new_n325_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT99), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n376_), .A2(new_n325_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n376_), .A2(new_n325_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(KEYINPUT4), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n430_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n434_), .A2(new_n435_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n430_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n429_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n436_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n428_), .B(new_n442_), .C1(new_n443_), .C2(new_n439_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n423_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n439_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT33), .B1(new_n448_), .B2(new_n429_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n348_), .B(KEYINPUT92), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n347_), .B1(new_n450_), .B2(new_n350_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT93), .B(new_n347_), .C1(new_n450_), .C2(new_n350_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n453_), .A2(new_n334_), .A3(new_n344_), .A4(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n339_), .B(KEYINPUT94), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n338_), .B1(new_n456_), .B2(G176gat), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n399_), .A2(new_n396_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n455_), .A2(new_n457_), .B1(new_n458_), .B2(new_n394_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n400_), .A2(new_n355_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT91), .Z(new_n464_));
  XOR2_X1   g263(.A(new_n464_), .B(KEYINPUT19), .Z(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT95), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT95), .ZN(new_n467_));
  INV_X1    g266(.A(new_n465_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n455_), .A2(new_n457_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n400_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT20), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n467_), .B(new_n468_), .C1(new_n471_), .C2(new_n460_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n400_), .A2(new_n355_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(KEYINPUT20), .C1(new_n469_), .C2(new_n400_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n474_), .A2(new_n468_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT97), .B(G8gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT98), .ZN(new_n484_));
  INV_X1    g283(.A(new_n482_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n466_), .A2(new_n472_), .A3(new_n485_), .A4(new_n475_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n483_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n476_), .A2(KEYINPUT98), .A3(new_n482_), .ZN(new_n488_));
  AOI211_X1 g287(.A(new_n445_), .B(new_n449_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n448_), .A2(new_n429_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n441_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(KEYINPUT32), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT101), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(new_n476_), .B2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n474_), .A2(new_n468_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n465_), .B2(new_n462_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n493_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n497_), .B(new_n498_), .C1(new_n476_), .C2(KEYINPUT101), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n492_), .B1(new_n495_), .B2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n362_), .B(new_n422_), .C1(new_n489_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT27), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n487_), .A2(new_n502_), .A3(new_n488_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n486_), .B(KEYINPUT27), .C1(new_n497_), .C2(new_n485_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n362_), .A2(new_n421_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n417_), .A2(new_n361_), .A3(new_n420_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n508_), .A3(new_n492_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n321_), .B1(new_n501_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n296_), .B(new_n241_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G231gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT16), .B(G183gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(G211gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(G127gat), .B(G155gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  OR3_X1    g318(.A1(new_n514_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(KEYINPUT17), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G134gat), .ZN(new_n525_));
  INV_X1    g324(.A(G162gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT75), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT72), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT34), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n307_), .A2(new_n308_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n538_), .A2(new_n243_), .B1(new_n534_), .B2(new_n533_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n234_), .A2(new_n288_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n537_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n536_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n539_), .A2(new_n536_), .A3(new_n535_), .A4(new_n540_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n530_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n527_), .B(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n543_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n546_), .B(new_n549_), .C1(new_n552_), .C2(new_n551_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n523_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT78), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n510_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n492_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n290_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT38), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n546_), .A2(new_n549_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(new_n523_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n510_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(G1gat), .B1(new_n564_), .B2(new_n492_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(G1324gat));
  INV_X1    g365(.A(KEYINPUT102), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT39), .ZN(new_n568_));
  OAI211_X1 g367(.A(G8gat), .B(new_n568_), .C1(new_n564_), .C2(new_n505_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(KEYINPUT39), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n505_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n558_), .A2(new_n291_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n570_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n571_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g375(.A(G15gat), .B1(new_n564_), .B2(new_n362_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT41), .Z(new_n578_));
  INV_X1    g377(.A(G15gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n362_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n558_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT103), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(G1326gat));
  OAI21_X1  g382(.A(G22gat), .B1(new_n564_), .B2(new_n422_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT42), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n422_), .A2(G22gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT104), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n558_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(G1327gat));
  AOI21_X1  g388(.A(new_n550_), .B1(new_n501_), .B2(new_n509_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n523_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n321_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(G29gat), .B1(new_n594_), .B2(new_n559_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT43), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n501_), .A2(new_n509_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n554_), .A2(new_n555_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n596_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  AOI211_X1 g399(.A(KEYINPUT43), .B(new_n598_), .C1(new_n501_), .C2(new_n509_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n592_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT44), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT44), .B(new_n592_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n604_), .A2(new_n559_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n595_), .B1(new_n606_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n572_), .A3(new_n605_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G36gat), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n593_), .A2(G36gat), .A3(new_n505_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT45), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT105), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(KEYINPUT46), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n609_), .B(new_n612_), .C1(new_n614_), .C2(KEYINPUT46), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1329gat));
  NAND4_X1  g417(.A1(new_n604_), .A2(G43gat), .A3(new_n361_), .A4(new_n605_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n282_), .B1(new_n593_), .B2(new_n362_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g421(.A1(new_n604_), .A2(new_n421_), .A3(new_n605_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G50gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n594_), .A2(new_n286_), .A3(new_n421_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT106), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT106), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n628_), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1331gat));
  INV_X1    g429(.A(new_n280_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n557_), .A2(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT107), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(KEYINPUT107), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n633_), .A2(new_n319_), .A3(new_n597_), .A4(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n492_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(G57gat), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n280_), .A2(new_n320_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n597_), .A2(new_n563_), .A3(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n492_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n637_), .B1(G57gat), .B2(new_n640_), .ZN(G1332gat));
  OAI21_X1  g440(.A(G64gat), .B1(new_n639_), .B2(new_n505_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT48), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n505_), .A2(G64gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n635_), .B2(new_n644_), .ZN(G1333gat));
  OR3_X1    g444(.A1(new_n635_), .A2(G71gat), .A3(new_n362_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G71gat), .B1(new_n639_), .B2(new_n362_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT108), .Z(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT49), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT49), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1334gat));
  OAI21_X1  g450(.A(G78gat), .B1(new_n639_), .B2(new_n422_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT50), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n422_), .A2(G78gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n635_), .B2(new_n654_), .ZN(G1335gat));
  NOR3_X1   g454(.A1(new_n280_), .A2(new_n320_), .A3(new_n591_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n590_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G85gat), .B1(new_n658_), .B2(new_n559_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n600_), .A2(new_n601_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n656_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n226_), .A2(new_n227_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n559_), .B1(new_n229_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT109), .Z(new_n665_));
  AOI21_X1  g464(.A(new_n659_), .B1(new_n662_), .B2(new_n665_), .ZN(G1336gat));
  NAND3_X1  g465(.A1(new_n662_), .A2(G92gat), .A3(new_n572_), .ZN(new_n667_));
  INV_X1    g466(.A(G92gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n668_), .B1(new_n657_), .B2(new_n505_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n667_), .A2(KEYINPUT110), .A3(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1337gat));
  OAI21_X1  g473(.A(G99gat), .B1(new_n661_), .B2(new_n362_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n658_), .A2(new_n222_), .A3(new_n361_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT51), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(KEYINPUT111), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n677_), .B(new_n679_), .ZN(G1338gat));
  OAI211_X1 g479(.A(new_n421_), .B(new_n656_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(G106gat), .A3(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n590_), .A2(new_n223_), .A3(new_n421_), .A4(new_n656_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT112), .ZN(new_n687_));
  INV_X1    g486(.A(new_n684_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n681_), .A2(G106gat), .A3(new_n688_), .A4(new_n682_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n687_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT53), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT53), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n685_), .A2(new_n692_), .A3(new_n687_), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1339gat));
  NOR2_X1   g493(.A1(new_n572_), .A2(new_n492_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n507_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT117), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT57), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n248_), .A2(new_n242_), .A3(new_n247_), .A4(new_n250_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n242_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n257_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(KEYINPUT55), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT55), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n701_), .A2(new_n704_), .A3(new_n257_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n272_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n319_), .B1(new_n706_), .B2(KEYINPUT114), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(KEYINPUT56), .ZN(new_n708_));
  INV_X1    g507(.A(new_n250_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n249_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n248_), .B1(new_n711_), .B2(new_n242_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n251_), .B1(new_n712_), .B2(new_n704_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n705_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT114), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT56), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .A4(new_n272_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n707_), .A2(new_n270_), .A3(new_n708_), .A4(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n306_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n303_), .A2(new_n304_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n301_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n315_), .A3(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n719_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n699_), .B1(new_n726_), .B2(new_n550_), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT57), .B(new_n562_), .C1(new_n719_), .C2(new_n725_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n724_), .A2(new_n270_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n715_), .A2(new_n717_), .A3(new_n272_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT115), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n270_), .A3(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n731_), .A2(new_n708_), .A3(new_n732_), .A4(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT58), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(KEYINPUT116), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(KEYINPUT116), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n598_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n698_), .B1(new_n729_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n735_), .A2(KEYINPUT116), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT58), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n735_), .A2(KEYINPUT116), .A3(new_n736_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n599_), .A3(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(KEYINPUT117), .C1(new_n727_), .C2(new_n728_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n523_), .A3(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n556_), .A2(new_n319_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT54), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n697_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G113gat), .B1(new_n749_), .B2(new_n320_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n697_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n729_), .A2(new_n739_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n591_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n748_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n751_), .B(new_n752_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT59), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n320_), .B(new_n756_), .C1(new_n749_), .C2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n750_), .B1(new_n759_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g559(.A(new_n324_), .B1(new_n280_), .B2(KEYINPUT60), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n749_), .B(new_n761_), .C1(KEYINPUT60), .C2(new_n324_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n631_), .B(new_n756_), .C1(new_n749_), .C2(new_n757_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(new_n324_), .ZN(G1341gat));
  INV_X1    g564(.A(G127gat), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n523_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n756_), .B(new_n767_), .C1(new_n749_), .C2(new_n757_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n749_), .A2(new_n591_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(G127gat), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT119), .ZN(G1342gat));
  AOI21_X1  g570(.A(G134gat), .B1(new_n749_), .B2(new_n562_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n772_), .A2(KEYINPUT120), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(KEYINPUT120), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n599_), .A2(G134gat), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n756_), .B(new_n775_), .C1(new_n749_), .C2(new_n757_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n773_), .A2(new_n774_), .A3(new_n776_), .ZN(G1343gat));
  AOI21_X1  g576(.A(new_n506_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n695_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n778_), .B2(new_n695_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n320_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT122), .B(G141gat), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n320_), .B(new_n784_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1344gat));
  OAI21_X1  g587(.A(new_n631_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G148gat), .ZN(new_n790_));
  INV_X1    g589(.A(G148gat), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n631_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1345gat));
  OAI21_X1  g592(.A(new_n591_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT61), .B(G155gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT123), .Z(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n796_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n591_), .B(new_n798_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1346gat));
  INV_X1    g599(.A(new_n782_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n526_), .B1(new_n801_), .B2(new_n780_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n562_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n599_), .A2(new_n802_), .B1(new_n803_), .B2(new_n526_), .ZN(G1347gat));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n505_), .A2(new_n559_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n580_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n422_), .B(new_n808_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n319_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n810_), .B2(new_n312_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT124), .B(G169gat), .C1(new_n809_), .C2(new_n319_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(KEYINPUT62), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT62), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n805_), .B(new_n814_), .C1(new_n810_), .C2(new_n312_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n810_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n813_), .B(new_n815_), .C1(new_n456_), .C2(new_n816_), .ZN(G1348gat));
  NAND2_X1  g616(.A1(new_n746_), .A2(new_n748_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n422_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT125), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n280_), .A2(new_n264_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT125), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n822_), .A3(new_n422_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n820_), .A2(new_n808_), .A3(new_n821_), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT126), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n264_), .B1(new_n809_), .B2(new_n280_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n822_), .B1(new_n818_), .B2(new_n422_), .ZN(new_n827_));
  AOI211_X1 g626(.A(KEYINPUT125), .B(new_n421_), .C1(new_n746_), .C2(new_n748_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT126), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n808_), .A4(new_n821_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n825_), .A2(new_n826_), .A3(new_n831_), .ZN(G1349gat));
  NAND2_X1  g631(.A1(new_n591_), .A2(new_n450_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n809_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n591_), .A3(new_n808_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n335_), .ZN(G1350gat));
  OR3_X1    g635(.A1(new_n809_), .A2(new_n350_), .A3(new_n550_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n809_), .A2(new_n598_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n336_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT127), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT127), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n837_), .B(new_n841_), .C1(new_n336_), .C2(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1351gat));
  NAND3_X1  g642(.A1(new_n778_), .A2(new_n320_), .A3(new_n806_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g644(.A1(new_n778_), .A2(new_n631_), .A3(new_n806_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g646(.A1(new_n778_), .A2(new_n591_), .A3(new_n806_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n849_));
  AND2_X1   g648(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n848_), .B2(new_n849_), .ZN(G1354gat));
  AND3_X1   g651(.A1(new_n778_), .A2(G218gat), .A3(new_n806_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n778_), .A2(new_n562_), .A3(new_n806_), .ZN(new_n854_));
  INV_X1    g653(.A(G218gat), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n853_), .A2(new_n599_), .B1(new_n854_), .B2(new_n855_), .ZN(G1355gat));
endmodule


