//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AND3_X1   g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(KEYINPUT85), .A3(new_n205_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G183gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT25), .B1(new_n218_), .B2(KEYINPUT84), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT84), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(G183gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(new_n203_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n223_), .A2(new_n227_), .B1(KEYINPUT24), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(KEYINPUT87), .A2(G176gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT87), .A2(G176gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT22), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n232_), .A2(new_n233_), .B1(new_n235_), .B2(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G169gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n237_), .A3(KEYINPUT22), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n229_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n208_), .A2(new_n240_), .A3(new_n209_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n217_), .A2(new_n231_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G204gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G197gat), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G204gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT96), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n245_), .B2(G204gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT21), .ZN(new_n250_));
  AND2_X1   g049(.A1(G211gat), .A2(G218gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G211gat), .A2(G218gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n247_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n255_), .A2(KEYINPUT21), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n244_), .A2(new_n246_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n257_), .A2(new_n255_), .A3(KEYINPUT21), .A4(new_n249_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n202_), .B1(new_n242_), .B2(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n254_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n219_), .A2(new_n222_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G169gat), .B(G176gat), .ZN(new_n263_));
  OAI22_X1  g062(.A1(new_n262_), .A2(new_n226_), .B1(new_n263_), .B2(new_n204_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n236_), .A2(new_n238_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n266_), .A2(new_n228_), .A3(new_n241_), .ZN(new_n267_));
  OAI211_X1 g066(.A(KEYINPUT100), .B(new_n261_), .C1(new_n265_), .C2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n260_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT20), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT101), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n237_), .A2(KEYINPUT22), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G169gat), .ZN(new_n277_));
  AND2_X1   g076(.A1(KEYINPUT87), .A2(G176gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(KEYINPUT87), .A2(G176gat), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n275_), .B(new_n277_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n228_), .A2(KEYINPUT99), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n228_), .A2(KEYINPUT99), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n280_), .A2(new_n241_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n285_));
  OAI22_X1  g084(.A1(new_n225_), .A2(new_n224_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n204_), .A2(KEYINPUT98), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT98), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT24), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n289_), .A3(new_n203_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n215_), .A3(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n263_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n283_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n274_), .B1(new_n261_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n293_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(new_n215_), .A3(new_n286_), .A4(new_n290_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n297_), .A2(new_n259_), .A3(KEYINPUT101), .A4(new_n283_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n273_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n269_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT102), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n261_), .A2(new_n294_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n242_), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT20), .B(new_n303_), .C1(new_n304_), .C2(new_n261_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n271_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n269_), .A2(new_n299_), .A3(KEYINPUT102), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT18), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(G64gat), .ZN(new_n311_));
  INV_X1    g110(.A(G92gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT103), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n302_), .A2(new_n306_), .A3(new_n307_), .A4(new_n313_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n302_), .A2(new_n307_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(KEYINPUT103), .A3(new_n306_), .A4(new_n313_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT104), .ZN(new_n322_));
  INV_X1    g121(.A(G155gat), .ZN(new_n323_));
  INV_X1    g122(.A(G162gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT92), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(G155gat), .A3(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT1), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT91), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G141gat), .B(G148gat), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337_));
  INV_X1    g136(.A(G141gat), .ZN(new_n338_));
  INV_X1    g137(.A(G148gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n331_), .A2(new_n345_), .A3(new_n328_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(KEYINPUT93), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT93), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n331_), .A2(new_n345_), .A3(new_n348_), .A4(new_n328_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n322_), .B(new_n336_), .C1(new_n347_), .C2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G120gat), .ZN(new_n352_));
  INV_X1    g151(.A(G127gat), .ZN(new_n353_));
  INV_X1    g152(.A(G134gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G127gat), .A2(G134gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT89), .ZN(new_n358_));
  INV_X1    g157(.A(G113gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT89), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n355_), .A2(new_n360_), .A3(new_n356_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n359_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n352_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(G120gat), .A3(new_n362_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n351_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n346_), .A2(KEYINPUT93), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n370_), .A2(new_n349_), .B1(new_n335_), .B2(new_n334_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n371_), .A2(new_n322_), .B1(new_n367_), .B2(new_n365_), .ZN(new_n372_));
  OR3_X1    g171(.A1(new_n369_), .A2(new_n372_), .A3(KEYINPUT107), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT105), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT107), .B1(new_n369_), .B2(new_n372_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G85gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT0), .ZN(new_n381_));
  INV_X1    g180(.A(G57gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT4), .B1(new_n369_), .B2(new_n372_), .ZN(new_n385_));
  OR3_X1    g184(.A1(new_n368_), .A2(KEYINPUT4), .A3(new_n371_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n374_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n378_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n376_), .A3(new_n386_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n374_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n383_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT106), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT33), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n321_), .A2(new_n388_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n305_), .A2(new_n271_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n269_), .B(KEYINPUT20), .C1(new_n261_), .C2(new_n294_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n271_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n313_), .A2(KEYINPUT32), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n400_), .B(new_n401_), .C1(new_n308_), .C2(KEYINPUT108), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT108), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n308_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n389_), .A2(new_n390_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n384_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n391_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n397_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT88), .B(KEYINPUT30), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n304_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n368_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n411_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n242_), .A2(new_n414_), .ZN(new_n415_));
  OR3_X1    g214(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n413_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G15gat), .B(G43gat), .Z(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n421_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n418_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430_));
  OAI211_X1 g229(.A(KEYINPUT95), .B(new_n261_), .C1(new_n371_), .C2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n430_), .B(new_n336_), .C1(new_n347_), .C2(new_n350_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT28), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT28), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n371_), .A2(new_n436_), .A3(new_n430_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n431_), .A2(new_n435_), .A3(new_n432_), .A4(new_n437_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G22gat), .B(G50gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT97), .B(new_n261_), .C1(new_n371_), .C2(new_n430_), .ZN(new_n445_));
  INV_X1    g244(.A(G228gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n451_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n445_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n443_), .A2(new_n444_), .A3(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n452_), .A2(new_n454_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n440_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n432_), .A2(new_n431_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n441_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n410_), .A2(new_n429_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n318_), .A2(new_n466_), .A3(new_n320_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT109), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n318_), .A2(KEYINPUT109), .A3(new_n466_), .A4(new_n320_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n418_), .B(new_n426_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n456_), .B2(new_n462_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n455_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n460_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n429_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n408_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n400_), .A2(new_n313_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(KEYINPUT27), .A3(new_n317_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n465_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G71gat), .B(G78gat), .Z(new_n482_));
  INV_X1    g281(.A(G64gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n382_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G57gat), .A2(G64gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT67), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n482_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n484_), .A2(new_n486_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(new_n485_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n489_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT10), .B(G99gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT65), .B(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(G92gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n312_), .A2(G85gat), .ZN(new_n512_));
  INV_X1    g311(.A(G85gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G92gat), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n504_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n502_), .A2(new_n505_), .A3(new_n511_), .A4(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  INV_X1    g317(.A(G99gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n501_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n508_), .A3(new_n521_), .A4(new_n509_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n512_), .A2(new_n514_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT8), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n521_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT66), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT66), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n520_), .A2(new_n528_), .A3(new_n521_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n527_), .A2(new_n511_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(KEYINPUT8), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n517_), .B(new_n525_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n498_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n499_), .A2(G106gat), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n534_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n524_), .B1(new_n535_), .B2(new_n505_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n527_), .A2(new_n511_), .A3(new_n529_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(KEYINPUT8), .A3(new_n523_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n496_), .A2(new_n536_), .A3(new_n497_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT64), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT68), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n533_), .A2(KEYINPUT12), .A3(new_n539_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n498_), .A2(new_n547_), .A3(new_n532_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n542_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(KEYINPUT68), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G120gat), .B(G148gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT5), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G176gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n243_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n545_), .A2(new_n550_), .A3(new_n551_), .A4(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT13), .Z(new_n561_));
  INV_X1    g360(.A(KEYINPUT83), .ZN(new_n562_));
  AND2_X1   g361(.A1(G29gat), .A2(G36gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(G29gat), .A2(G36gat), .ZN(new_n564_));
  OAI21_X1  g363(.A(G43gat), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(G29gat), .ZN(new_n566_));
  INV_X1    g365(.A(G36gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(G43gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G29gat), .A2(G36gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(G50gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(new_n571_), .A3(G50gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G8gat), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT74), .B(G8gat), .ZN(new_n581_));
  INV_X1    g380(.A(G1gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT14), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n580_), .A2(new_n585_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n577_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n578_), .B(KEYINPUT75), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n580_), .A2(new_n585_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n576_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT79), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT15), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n565_), .A2(new_n571_), .A3(G50gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(G50gat), .B1(new_n565_), .B2(new_n571_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n574_), .A2(KEYINPUT15), .A3(new_n575_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n590_), .A2(new_n591_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n588_), .B(new_n594_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT79), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n593_), .A2(new_n607_), .A3(new_n595_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n597_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT82), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT80), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(G169gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G197gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n613_), .B(new_n237_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n245_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(KEYINPUT81), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT81), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n609_), .A2(new_n610_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n610_), .B1(new_n609_), .B2(new_n622_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n597_), .A2(new_n606_), .A3(new_n608_), .A4(new_n618_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n562_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n609_), .A2(new_n622_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT82), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n609_), .A2(new_n622_), .A3(new_n610_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n629_), .A2(new_n562_), .A3(new_n626_), .A4(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n561_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n481_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT69), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT34), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT35), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n536_), .A2(new_n577_), .A3(KEYINPUT70), .A4(new_n538_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT70), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n532_), .B2(new_n603_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n532_), .A2(new_n576_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n640_), .B(new_n641_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n638_), .A2(new_n639_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n536_), .A2(new_n538_), .B1(new_n602_), .B2(new_n601_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n648_), .A2(new_n642_), .B1(new_n532_), .B2(new_n576_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n646_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n640_), .A4(new_n641_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT72), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G190gat), .B(G218gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(G134gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(new_n324_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT36), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT72), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n647_), .A2(new_n651_), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT36), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n652_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT71), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n657_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n657_), .A2(new_n667_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n652_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT37), .B1(new_n670_), .B2(new_n663_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n498_), .B(new_n605_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(G231gat), .A2(G233gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT76), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n674_), .B(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n678_));
  XNOR2_X1  g477(.A(G127gat), .B(G155gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(G183gat), .B(G211gat), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n680_), .B(new_n681_), .Z(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT78), .B1(new_n683_), .B2(KEYINPUT17), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n677_), .A2(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n683_), .A2(KEYINPUT17), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n677_), .A2(new_n685_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n673_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n635_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n582_), .A3(new_n408_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT38), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT110), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT110), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n660_), .A2(new_n664_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n689_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n635_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n582_), .B1(new_n701_), .B2(new_n408_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n696_), .A2(new_n697_), .A3(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n694_), .B2(new_n693_), .ZN(G1324gat));
  INV_X1    g503(.A(new_n479_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n692_), .A2(new_n581_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n701_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G8gat), .B1(new_n709_), .B2(new_n706_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT39), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT39), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT40), .B(new_n708_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1325gat));
  OAI21_X1  g516(.A(G15gat), .B1(new_n709_), .B2(new_n429_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT41), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n691_), .A2(G15gat), .A3(new_n429_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1326gat));
  NOR2_X1   g520(.A1(new_n464_), .A2(G22gat), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT111), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n692_), .A2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G22gat), .B1(new_n709_), .B2(new_n464_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(KEYINPUT42), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(KEYINPUT42), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(new_n724_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1327gat));
  NAND3_X1  g531(.A1(new_n666_), .A2(new_n671_), .A3(KEYINPUT113), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT43), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n463_), .B1(new_n397_), .B2(new_n409_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n429_), .A2(new_n735_), .B1(new_n706_), .B2(new_n477_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n736_), .B2(new_n672_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n734_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n481_), .A2(new_n673_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n689_), .A3(new_n634_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n740_), .A2(KEYINPUT44), .A3(new_n689_), .A4(new_n634_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n408_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G29gat), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n689_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(new_n698_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n635_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n566_), .A3(new_n408_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n751_), .ZN(G1328gat));
  OAI21_X1  g551(.A(G36gat), .B1(new_n745_), .B2(new_n706_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n567_), .A3(new_n707_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT45), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n753_), .B(new_n755_), .C1(KEYINPUT114), .C2(KEYINPUT46), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1329gat));
  OAI21_X1  g559(.A(G43gat), .B1(new_n745_), .B2(new_n429_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n750_), .A2(new_n569_), .A3(new_n472_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(KEYINPUT47), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1330gat));
  OAI21_X1  g566(.A(G50gat), .B1(new_n745_), .B2(new_n464_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n750_), .A2(new_n573_), .A3(new_n463_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1331gat));
  INV_X1    g569(.A(new_n633_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n736_), .A2(new_n771_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT115), .Z(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(new_n561_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n408_), .A3(new_n690_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n772_), .A2(new_n561_), .A3(new_n700_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n746_), .A2(new_n382_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n775_), .A2(new_n382_), .B1(new_n776_), .B2(new_n777_), .ZN(G1332gat));
  INV_X1    g577(.A(new_n776_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G64gat), .B1(new_n779_), .B2(new_n706_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT48), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT48), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n690_), .A3(new_n561_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n707_), .A2(new_n483_), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n781_), .A2(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI221_X1 g586(.A(KEYINPUT116), .B1(new_n783_), .B2(new_n784_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1333gat));
  INV_X1    g588(.A(G71gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n776_), .B2(new_n472_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT49), .Z(new_n792_));
  NAND2_X1  g591(.A1(new_n472_), .A2(new_n790_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n783_), .B2(new_n793_), .ZN(G1334gat));
  INV_X1    g593(.A(G78gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n776_), .B2(new_n463_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT50), .Z(new_n797_));
  NAND2_X1  g596(.A1(new_n463_), .A2(new_n795_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n783_), .B2(new_n798_), .ZN(G1335gat));
  NAND3_X1  g598(.A1(new_n773_), .A2(new_n561_), .A3(new_n749_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G85gat), .B1(new_n801_), .B2(new_n408_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n560_), .B(KEYINPUT13), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n771_), .A2(new_n803_), .A3(new_n748_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n740_), .A2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n408_), .A2(new_n503_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(G1336gat));
  AOI21_X1  g606(.A(G92gat), .B1(new_n801_), .B2(new_n707_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n706_), .A2(new_n312_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n805_), .B2(new_n809_), .ZN(G1337gat));
  INV_X1    g609(.A(new_n805_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G99gat), .B1(new_n811_), .B2(new_n429_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n472_), .A2(new_n500_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n800_), .B2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g614(.A(new_n738_), .B1(new_n481_), .B2(new_n673_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n672_), .B(new_n734_), .C1(new_n465_), .C2(new_n480_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n463_), .B(new_n804_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT117), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n740_), .A2(new_n820_), .A3(new_n463_), .A4(new_n804_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(G106gat), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT52), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n819_), .A2(new_n824_), .A3(new_n821_), .A4(G106gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n464_), .A2(G106gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n801_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT53), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1339gat));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n543_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n546_), .A2(new_n543_), .A3(new_n548_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT55), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n838_), .B(new_n556_), .C1(new_n840_), .C2(new_n836_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n550_), .A2(KEYINPUT55), .A3(new_n839_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(KEYINPUT56), .A3(new_n556_), .A4(new_n838_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n845_), .A3(KEYINPUT120), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(new_n559_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n845_), .A2(KEYINPUT120), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n629_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT83), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n850_), .B2(new_n631_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n593_), .A2(new_n594_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n588_), .B(new_n595_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n852_), .A2(new_n615_), .A3(new_n853_), .A4(new_n617_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n626_), .A2(new_n854_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n847_), .A2(new_n851_), .B1(new_n560_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n835_), .B1(new_n856_), .B2(new_n699_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n560_), .A2(new_n855_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n848_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n846_), .A2(new_n559_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(KEYINPUT57), .A3(new_n698_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n843_), .A2(new_n845_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n559_), .A3(new_n855_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n866_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n673_), .A3(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n857_), .A2(new_n863_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n689_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n690_), .A2(new_n633_), .A3(new_n803_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT54), .Z(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n690_), .A2(new_n633_), .A3(new_n803_), .A4(new_n874_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n871_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n707_), .A2(new_n746_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n473_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT122), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n880_), .A2(KEYINPUT123), .A3(new_n881_), .A4(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n878_), .B1(new_n870_), .B2(new_n689_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT59), .B1(new_n887_), .B2(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n633_), .A2(new_n359_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT59), .B1(new_n871_), .B2(new_n879_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT123), .B1(new_n892_), .B2(new_n885_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n889_), .A2(new_n891_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n884_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n880_), .A2(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(KEYINPUT121), .B(new_n359_), .C1(new_n896_), .C2(new_n633_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n887_), .A2(new_n633_), .A3(new_n884_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(G113gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n834_), .B1(new_n894_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n892_), .A2(new_n885_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n905_), .A2(new_n890_), .A3(new_n888_), .A4(new_n886_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n906_), .A2(KEYINPUT124), .A3(new_n900_), .A4(new_n897_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n907_), .ZN(G1340gat));
  AOI21_X1  g707(.A(KEYINPUT60), .B1(new_n561_), .B2(new_n352_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n887_), .A2(new_n884_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n889_), .A2(new_n893_), .A3(new_n910_), .A4(new_n803_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n352_), .ZN(G1341gat));
  INV_X1    g713(.A(new_n896_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G127gat), .B1(new_n915_), .B2(new_n748_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n889_), .A2(new_n893_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n689_), .A2(new_n353_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1342gat));
  AOI21_X1  g718(.A(G134gat), .B1(new_n915_), .B2(new_n699_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n672_), .A2(new_n354_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n917_), .B2(new_n921_), .ZN(G1343gat));
  NOR2_X1   g721(.A1(new_n887_), .A2(new_n476_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n882_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n633_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n338_), .ZN(G1344gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n803_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n339_), .ZN(G1345gat));
  NOR2_X1   g727(.A1(new_n924_), .A2(new_n689_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT61), .B(G155gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  NOR3_X1   g730(.A1(new_n924_), .A2(new_n324_), .A3(new_n672_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n924_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n699_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n324_), .B2(new_n934_), .ZN(G1347gat));
  XOR2_X1   g734(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n887_), .A2(new_n473_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n938_), .A2(new_n746_), .A3(new_n707_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n633_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n937_), .B1(new_n940_), .B2(new_n237_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n940_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n942_));
  OAI211_X1 g741(.A(G169gat), .B(new_n936_), .C1(new_n939_), .C2(new_n633_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(G1348gat));
  NAND4_X1  g743(.A1(new_n938_), .A2(new_n746_), .A3(new_n561_), .A4(new_n707_), .ZN(new_n945_));
  INV_X1    g744(.A(G176gat), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n232_), .A2(new_n233_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n945_), .ZN(G1349gat));
  NOR2_X1   g748(.A1(new_n939_), .A2(new_n689_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(new_n285_), .B2(new_n284_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n951_), .B1(new_n218_), .B2(new_n950_), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n939_), .B2(new_n672_), .ZN(new_n953_));
  OR2_X1    g752(.A1(new_n939_), .A2(new_n226_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n698_), .ZN(G1351gat));
  NOR2_X1   g754(.A1(new_n887_), .A2(new_n706_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n476_), .A2(new_n408_), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT126), .Z(new_n958_));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n633_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(new_n245_), .ZN(G1352gat));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n803_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(new_n243_), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n956_), .A2(new_n748_), .A3(new_n958_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  AND2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n964_), .A2(new_n965_), .A3(new_n966_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(new_n964_), .B2(new_n965_), .ZN(G1354gat));
  INV_X1    g767(.A(G218gat), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n969_), .B1(new_n959_), .B2(new_n698_), .ZN(new_n970_));
  NAND4_X1  g769(.A1(new_n956_), .A2(G218gat), .A3(new_n673_), .A4(new_n958_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(KEYINPUT127), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n970_), .A2(new_n974_), .A3(new_n971_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n975_), .ZN(G1355gat));
endmodule


