//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n205_), .A2(KEYINPUT24), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT23), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n209_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT22), .B(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n214_), .A3(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n207_), .B(new_n219_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n216_), .A2(KEYINPUT30), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT30), .B1(new_n216_), .B2(new_n225_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT77), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT76), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G71gat), .B(G99gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G15gat), .B(G43gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n229_), .A2(new_n230_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n236_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(new_n228_), .C1(new_n227_), .C2(new_n226_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT31), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT31), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n237_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT78), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G127gat), .B(G134gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT78), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n248_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n250_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n249_), .A2(KEYINPUT79), .A3(new_n251_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n247_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n243_), .A2(new_n258_), .A3(new_n257_), .A4(new_n246_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT81), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(KEYINPUT82), .A3(new_n266_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT3), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT2), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n271_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n265_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n266_), .B(KEYINPUT1), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n273_), .B(new_n277_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT29), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT84), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G197gat), .A2(G204gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT83), .B(G204gat), .Z(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(G197gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(KEYINPUT21), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(G197gat), .B2(G204gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n287_), .B2(G197gat), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n292_), .B(new_n283_), .C1(new_n288_), .C2(KEYINPUT21), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT86), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT86), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n282_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G228gat), .A3(G233gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G228gat), .A2(G233gat), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n282_), .A2(KEYINPUT85), .A3(new_n294_), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n294_), .A2(new_n300_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n302_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n299_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G78gat), .B(G106gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n276_), .A2(new_n303_), .A3(new_n280_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G22gat), .B(G50gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT28), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n313_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n299_), .A2(new_n307_), .A3(KEYINPUT87), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT87), .B1(new_n299_), .B2(new_n307_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n310_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n308_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n299_), .A2(new_n307_), .A3(KEYINPUT87), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(KEYINPUT88), .A3(new_n310_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n318_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n308_), .A2(new_n310_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n317_), .B1(new_n312_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n262_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n318_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT88), .B1(new_n327_), .B2(new_n310_), .ZN(new_n334_));
  AOI211_X1 g133(.A(new_n322_), .B(new_n311_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n260_), .A2(new_n261_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n332_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n223_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n209_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n207_), .A2(KEYINPUT89), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n207_), .A2(KEYINPUT89), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n343_), .A2(new_n219_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n294_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n216_), .A2(new_n225_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n348_), .B(KEYINPUT20), .C1(new_n294_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT90), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G64gat), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(G92gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(G92gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n347_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n289_), .A2(new_n293_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n352_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n349_), .A2(new_n294_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n364_), .A2(KEYINPUT20), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n354_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n353_), .A2(KEYINPUT90), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n367_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n360_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT27), .B1(new_n368_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n252_), .A2(new_n255_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n281_), .A2(new_n376_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n257_), .A2(new_n258_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n379_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n375_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n377_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n259_), .A2(new_n281_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT4), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n388_), .A2(KEYINPUT91), .A3(new_n383_), .A4(new_n381_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n382_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n385_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT0), .ZN(new_n393_));
  INV_X1    g192(.A(G57gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n385_), .A2(new_n389_), .A3(new_n399_), .A4(new_n390_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n360_), .B(KEYINPUT95), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n363_), .A2(new_n296_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n297_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n362_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT20), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n406_), .A2(KEYINPUT93), .B1(new_n294_), .B2(new_n349_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT93), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n408_), .A3(KEYINPUT20), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n365_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n410_), .A2(KEYINPUT94), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n350_), .A2(new_n352_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n410_), .B2(KEYINPUT94), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n402_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n368_), .A2(KEYINPUT27), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n374_), .B(new_n401_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n372_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n398_), .A2(new_n400_), .B1(new_n420_), .B2(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n400_), .B(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n388_), .A2(new_n382_), .A3(new_n381_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n386_), .A2(new_n387_), .A3(new_n383_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n397_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n368_), .A2(new_n373_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n423_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n400_), .B(KEYINPUT33), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n368_), .A2(new_n373_), .A3(new_n428_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT92), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n329_), .A2(new_n338_), .A3(new_n331_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n340_), .A2(new_n416_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G229gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G29gat), .B(G36gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(KEYINPUT70), .ZN(new_n441_));
  INV_X1    g240(.A(G36gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G29gat), .ZN(new_n443_));
  INV_X1    g242(.A(G29gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G36gat), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n443_), .A2(new_n445_), .A3(KEYINPUT70), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n441_), .A2(new_n446_), .A3(G43gat), .ZN(new_n447_));
  INV_X1    g246(.A(G43gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n445_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT70), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n440_), .A2(KEYINPUT70), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n439_), .B1(new_n447_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  INV_X1    g254(.A(G1gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(G43gat), .B1(new_n441_), .B2(new_n446_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n451_), .A2(new_n452_), .A3(new_n448_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(G50gat), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n454_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(new_n454_), .B2(new_n465_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n438_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n454_), .A2(new_n465_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n454_), .A2(KEYINPUT15), .A3(new_n465_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n462_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n466_), .A2(new_n437_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G113gat), .B(G141gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G169gat), .ZN(new_n478_));
  INV_X1    g277(.A(G197gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n469_), .B(new_n480_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G232gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT34), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT10), .ZN(new_n489_));
  INV_X1    g288(.A(G99gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT64), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(KEYINPUT64), .A3(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(G106gat), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G92gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n396_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(KEYINPUT9), .A3(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT68), .B1(new_n496_), .B2(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n499_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n491_), .A2(KEYINPUT64), .A3(new_n492_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(new_n493_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n507_), .B(new_n508_), .C1(new_n510_), .C2(G106gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT66), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521_));
  NOR4_X1   g320(.A1(new_n521_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT65), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n520_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n501_), .B(new_n502_), .C1(KEYINPUT66), .C2(new_n512_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n514_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n521_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(KEYINPUT65), .A3(new_n524_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n530_), .A2(new_n499_), .A3(new_n519_), .A4(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n527_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n513_), .A3(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n506_), .A2(new_n511_), .A3(new_n528_), .A4(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n473_), .B2(new_n472_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n507_), .B1(new_n510_), .B2(G106gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n528_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n470_), .A2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT35), .B(new_n488_), .C1(new_n537_), .C2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n472_), .A2(new_n473_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n535_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n488_), .A2(KEYINPUT35), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n488_), .A2(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n540_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n541_), .A2(new_n545_), .A3(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n544_), .B(KEYINPUT36), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n541_), .B2(new_n552_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n486_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n552_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n549_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n554_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n541_), .A2(new_n545_), .A3(new_n552_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(KEYINPUT37), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  INV_X1    g363(.A(G64gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G57gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n394_), .A2(G64gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT11), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n567_), .A3(KEYINPUT11), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(KEYINPUT11), .A3(new_n566_), .A4(new_n567_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT67), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(KEYINPUT67), .A3(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n539_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n581_), .A2(new_n582_), .B1(new_n535_), .B2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n532_), .A2(new_n513_), .A3(new_n533_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n513_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n587_), .A2(new_n579_), .A3(new_n578_), .A4(new_n538_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT69), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(KEYINPUT69), .B(new_n589_), .C1(new_n580_), .C2(new_n539_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n584_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n589_), .B1(new_n588_), .B2(new_n581_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G120gat), .B(G148gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G204gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT5), .B(G176gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  NAND3_X1  g398(.A1(new_n593_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n564_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(KEYINPUT13), .A3(new_n600_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT16), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(G183gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n608_), .B(new_n210_), .ZN(new_n611_));
  INV_X1    g410(.A(G211gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT17), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT71), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n461_), .B(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n618_), .A2(new_n580_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n610_), .A2(new_n613_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n580_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n615_), .A2(new_n619_), .A3(new_n621_), .A4(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n576_), .B(KEYINPUT72), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n624_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(KEYINPUT17), .A3(new_n614_), .A4(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n623_), .A2(KEYINPUT73), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT73), .B1(new_n623_), .B2(new_n627_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n563_), .A2(new_n606_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT74), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  NOR4_X1   g434(.A1(new_n436_), .A2(new_n485_), .A3(new_n634_), .A4(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n401_), .B(KEYINPUT96), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n456_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT97), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n340_), .A2(new_n416_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n434_), .A2(new_n435_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n606_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n484_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n553_), .A2(new_n556_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT98), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n623_), .A2(new_n627_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n645_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n643_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n401_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n640_), .A2(new_n653_), .ZN(G1324gat));
  AOI21_X1  g453(.A(new_n374_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n457_), .B1(new_n650_), .B2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT39), .Z(new_n658_));
  NAND3_X1  g457(.A1(new_n636_), .A2(new_n457_), .A3(new_n656_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(G1325gat));
  INV_X1    g461(.A(G15gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n650_), .B2(new_n338_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT41), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n636_), .A2(new_n663_), .A3(new_n338_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT99), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n329_), .A2(new_n331_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(G22gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT100), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n636_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G22gat), .B1(new_n651_), .B2(new_n669_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(KEYINPUT42), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(KEYINPUT42), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(G1327gat));
  INV_X1    g475(.A(new_n646_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n436_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n645_), .A2(new_n630_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n401_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n643_), .B2(new_n563_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n563_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT43), .B(new_n685_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n679_), .C1(new_n684_), .C2(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(G29gat), .A3(new_n637_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n679_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n682_), .B1(new_n688_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(new_n679_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n436_), .B2(new_n685_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n643_), .A2(new_n683_), .A3(new_n563_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n655_), .B1(new_n696_), .B2(KEYINPUT44), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n442_), .B1(new_n697_), .B2(new_n691_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n656_), .A2(KEYINPUT101), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n656_), .A2(KEYINPUT101), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n442_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n680_), .A2(new_n699_), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n699_), .B1(new_n680_), .B2(new_n703_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n698_), .A2(new_n706_), .B1(KEYINPUT102), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(KEYINPUT102), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1329gat));
  OAI21_X1  g509(.A(new_n448_), .B1(new_n680_), .B2(new_n262_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT103), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n696_), .A2(KEYINPUT44), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n687_), .A2(G43gat), .A3(new_n338_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g515(.A(new_n669_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n687_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT104), .B1(new_n718_), .B2(new_n713_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n691_), .A2(new_n720_), .A3(new_n717_), .A4(new_n687_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n721_), .A3(G50gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n681_), .A2(new_n439_), .A3(new_n717_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT105), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n644_), .A2(new_n484_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n643_), .A2(new_n630_), .A3(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n563_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n637_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n730_), .A2(new_n647_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT106), .B(G57gat), .Z(new_n734_));
  NOR2_X1   g533(.A1(new_n652_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n732_), .B1(new_n733_), .B2(new_n735_), .ZN(G1332gat));
  AOI21_X1  g535(.A(new_n565_), .B1(new_n733_), .B2(new_n702_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT48), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n731_), .A2(new_n565_), .A3(new_n702_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n733_), .B2(new_n338_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT49), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n731_), .A2(new_n741_), .A3(new_n338_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT107), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(new_n747_), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1334gat));
  INV_X1    g548(.A(G78gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n731_), .A2(new_n750_), .A3(new_n717_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n733_), .A2(new_n717_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G78gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n754_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n751_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT109), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n729_), .A2(new_n631_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n678_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n396_), .A3(new_n637_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n760_), .A2(KEYINPUT110), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(KEYINPUT110), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n694_), .A2(new_n695_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(new_n401_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n767_), .B2(new_n396_), .ZN(G1336gat));
  OAI21_X1  g567(.A(new_n500_), .B1(new_n761_), .B2(new_n655_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT111), .Z(new_n770_));
  INV_X1    g569(.A(new_n702_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n500_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n766_), .B2(new_n772_), .ZN(G1337gat));
  AND2_X1   g572(.A1(new_n766_), .A2(new_n338_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n338_), .B1(new_n509_), .B2(new_n493_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n774_), .A2(new_n490_), .B1(new_n761_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT112), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n776_), .B(new_n778_), .ZN(G1338gat));
  INV_X1    g578(.A(G106gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n762_), .A2(new_n780_), .A3(new_n717_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n766_), .A2(new_n717_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G106gat), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT52), .B(new_n780_), .C1(new_n766_), .C2(new_n717_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT53), .ZN(G1339gat));
  XOR2_X1   g586(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n788_));
  OAI21_X1  g587(.A(new_n437_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n466_), .A2(new_n438_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n789_), .B(new_n481_), .C1(new_n474_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n483_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n483_), .A3(KEYINPUT116), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n604_), .A2(new_n600_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT55), .B(new_n584_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n589_), .B1(new_n580_), .B2(new_n539_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT69), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n591_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n803_), .B2(new_n584_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n589_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n799_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n797_), .B1(new_n806_), .B2(new_n599_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n599_), .A2(new_n797_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n806_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n593_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n805_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n798_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(KEYINPUT115), .A3(new_n809_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n807_), .A2(new_n811_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n484_), .A2(new_n600_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT114), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n484_), .A2(new_n820_), .A3(new_n600_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n796_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n788_), .B1(new_n823_), .B2(new_n646_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n821_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n599_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT115), .B1(new_n815_), .B2(new_n809_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n825_), .B1(new_n829_), .B2(new_n816_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT57), .B(new_n677_), .C1(new_n830_), .C2(new_n796_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT58), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n804_), .A2(new_n805_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n599_), .B1(new_n836_), .B2(new_n798_), .ZN(new_n837_));
  OAI22_X1  g636(.A1(new_n837_), .A2(KEYINPUT56), .B1(new_n806_), .B2(new_n810_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n601_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n835_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n810_), .B1(new_n836_), .B2(new_n798_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n839_), .B(new_n835_), .C1(new_n827_), .C2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n563_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n832_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n839_), .B1(new_n827_), .B2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n834_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(KEYINPUT119), .A3(new_n563_), .A4(new_n842_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n824_), .A2(new_n831_), .A3(new_n844_), .A4(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n648_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n557_), .A2(new_n630_), .A3(new_n562_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n850_), .A2(new_n644_), .A3(new_n851_), .A4(new_n485_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT113), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n644_), .A3(new_n485_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT54), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n852_), .A2(KEYINPUT113), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n849_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n339_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n655_), .A3(new_n637_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(G113gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n484_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n824_), .B(new_n831_), .C1(new_n840_), .C2(new_n843_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n631_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n858_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n862_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT120), .B1(new_n863_), .B2(KEYINPUT59), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n848_), .A2(new_n648_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n873_), .C2(new_n861_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n871_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT122), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n869_), .A2(new_n862_), .A3(new_n870_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT59), .B1(new_n873_), .B2(new_n861_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n878_), .B1(new_n881_), .B2(new_n874_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n485_), .B1(new_n877_), .B2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n866_), .B1(new_n885_), .B2(new_n865_), .ZN(G1340gat));
  OAI21_X1  g685(.A(G120gat), .B1(new_n876_), .B2(new_n644_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n644_), .A2(G120gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(KEYINPUT60), .ZN(new_n890_));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(KEYINPUT60), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n864_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n887_), .A2(new_n888_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n882_), .B2(new_n606_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n893_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT123), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(G1341gat));
  INV_X1    g697(.A(G127gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n864_), .A2(new_n899_), .A3(new_n630_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n648_), .B1(new_n877_), .B2(new_n884_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1342gat));
  AOI21_X1  g701(.A(G134gat), .B1(new_n864_), .B2(new_n647_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n877_), .A2(new_n884_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n563_), .A2(G134gat), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT124), .Z(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n904_), .B2(new_n906_), .ZN(G1343gat));
  NOR2_X1   g706(.A1(new_n873_), .A2(new_n332_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n637_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n702_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n484_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n606_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g715(.A1(new_n911_), .A2(new_n631_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT61), .B(G155gat), .Z(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n911_), .B2(new_n685_), .ZN(new_n920_));
  INV_X1    g719(.A(G162gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n647_), .A2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n911_), .B2(new_n922_), .ZN(G1347gat));
  NAND3_X1  g722(.A1(new_n702_), .A2(new_n338_), .A3(new_n909_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n717_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n869_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G169gat), .B1(new_n926_), .B2(new_n485_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT62), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n484_), .A2(new_n217_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT125), .Z(new_n930_));
  OAI21_X1  g729(.A(new_n928_), .B1(new_n926_), .B2(new_n930_), .ZN(G1348gat));
  INV_X1    g730(.A(new_n926_), .ZN(new_n932_));
  AOI21_X1  g731(.A(G176gat), .B1(new_n932_), .B2(new_n606_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n873_), .A2(new_n717_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n924_), .A2(new_n218_), .A3(new_n644_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(G1349gat));
  NOR3_X1   g735(.A1(new_n926_), .A2(new_n202_), .A3(new_n648_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n924_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n934_), .A2(new_n630_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n210_), .B2(new_n939_), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n926_), .B2(new_n685_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n647_), .A2(new_n203_), .ZN(new_n942_));
  XOR2_X1   g741(.A(new_n942_), .B(KEYINPUT126), .Z(new_n943_));
  OAI21_X1  g742(.A(new_n941_), .B1(new_n926_), .B2(new_n943_), .ZN(G1351gat));
  NOR2_X1   g743(.A1(new_n771_), .A2(new_n401_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n908_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n485_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n479_), .ZN(G1352gat));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n644_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(G204gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n950_), .B1(new_n287_), .B2(new_n949_), .ZN(G1353gat));
  INV_X1    g750(.A(new_n946_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n648_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT127), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n954_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n955_), .B(new_n956_), .Z(G1354gat));
  OAI21_X1  g756(.A(G218gat), .B1(new_n946_), .B2(new_n685_), .ZN(new_n958_));
  INV_X1    g757(.A(G218gat), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n647_), .A2(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n958_), .B1(new_n946_), .B2(new_n960_), .ZN(G1355gat));
endmodule


