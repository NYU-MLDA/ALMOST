//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203_));
  OR2_X1    g002(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT26), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT25), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n209_), .B(new_n211_), .C1(KEYINPUT26), .C2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n203_), .B1(new_n207_), .B2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n209_), .A2(new_n211_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n212_), .A2(KEYINPUT26), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n215_), .A2(new_n206_), .A3(KEYINPUT76), .A4(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224_));
  INV_X1    g023(.A(new_n222_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n219_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(KEYINPUT23), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n223_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n218_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n204_), .A2(new_n208_), .A3(new_n205_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n227_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(new_n230_), .C2(KEYINPUT78), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT22), .B(G169gat), .Z(new_n236_));
  OAI21_X1  g035(.A(new_n221_), .B1(new_n236_), .B2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT86), .B(G204gat), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G218gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G211gat), .ZN(new_n247_));
  INV_X1    g046(.A(G211gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G218gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT21), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT88), .B1(new_n245_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G204gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT86), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT86), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G204gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n244_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n258_), .A2(new_n259_), .A3(new_n261_), .A4(new_n242_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n252_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n260_), .B1(new_n257_), .B2(new_n241_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n256_), .A3(new_n244_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n260_), .B1(G197gat), .B2(G204gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n250_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n264_), .A2(KEYINPUT87), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT87), .B1(new_n264_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n263_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT20), .B1(new_n240_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(G190gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n215_), .A2(new_n272_), .ZN(new_n273_));
  OR3_X1    g072(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n223_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n234_), .B1(new_n230_), .B2(KEYINPUT78), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n228_), .A2(new_n229_), .B1(new_n208_), .B2(new_n212_), .ZN(new_n277_));
  OAI22_X1  g076(.A1(new_n275_), .A2(new_n276_), .B1(new_n237_), .B2(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT19), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n271_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT20), .B1(new_n270_), .B2(new_n278_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT94), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n240_), .A2(new_n270_), .ZN(new_n286_));
  OAI211_X1 g085(.A(KEYINPUT94), .B(KEYINPUT20), .C1(new_n270_), .C2(new_n278_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n288_), .B2(new_n281_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G64gat), .B(G92gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(G8gat), .B(G36gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT95), .B1(new_n289_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n281_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n286_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(new_n283_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT90), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n301_), .B(new_n281_), .C1(new_n271_), .C2(new_n279_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n264_), .A2(new_n267_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n264_), .A2(KEYINPUT87), .A3(new_n267_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n306_), .A2(new_n307_), .B1(new_n252_), .B2(new_n262_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n218_), .A2(new_n231_), .B1(new_n238_), .B2(new_n235_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n270_), .A2(new_n278_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT20), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n301_), .B1(new_n312_), .B2(new_n281_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n295_), .B(new_n300_), .C1(new_n303_), .C2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n283_), .A2(new_n284_), .B1(new_n240_), .B2(new_n270_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n297_), .B1(new_n316_), .B2(new_n287_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n315_), .B(new_n294_), .C1(new_n317_), .C2(new_n282_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n296_), .A2(KEYINPUT27), .A3(new_n314_), .A4(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n300_), .B1(new_n303_), .B2(new_n313_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n294_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT27), .B1(new_n321_), .B2(new_n314_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT27), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n281_), .B1(new_n271_), .B2(new_n279_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT90), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n302_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n295_), .B1(new_n328_), .B2(new_n300_), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n294_), .B(new_n299_), .C1(new_n327_), .C2(new_n302_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n325_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(KEYINPUT96), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n202_), .B1(new_n324_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G120gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n335_), .A2(new_n336_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n338_), .A2(G113gat), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G113gat), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n335_), .A2(new_n336_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n337_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n334_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(G113gat), .B1(new_n338_), .B2(new_n339_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n341_), .A3(new_n337_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(G120gat), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT31), .B1(new_n344_), .B2(new_n347_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT83), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n309_), .B(KEYINPUT30), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n354_), .A2(KEYINPUT80), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(KEYINPUT80), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G227gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT79), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G15gat), .B(G43gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(new_n356_), .A3(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(new_n354_), .A2(KEYINPUT80), .A3(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n353_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n364_), .A3(KEYINPUT81), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n367_), .A2(new_n368_), .B1(new_n352_), .B2(new_n365_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT84), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT3), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT2), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n374_), .B(new_n375_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n375_), .B(KEYINPUT1), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n374_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n376_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n379_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n372_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n371_), .B1(new_n389_), .B2(new_n308_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n374_), .A2(new_n375_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n377_), .A2(new_n380_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT85), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n393_), .B2(new_n381_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n388_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n270_), .B(new_n370_), .C1(new_n396_), .C2(new_n372_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n390_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n396_), .A2(new_n372_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G22gat), .B(G50gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT28), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n403_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n390_), .A2(new_n397_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n398_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n400_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n409_), .A2(KEYINPUT89), .A3(new_n400_), .A4(new_n406_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT0), .ZN(new_n416_));
  INV_X1    g215(.A(G57gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G85gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n384_), .A2(new_n388_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n348_), .A3(KEYINPUT92), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n396_), .A2(new_n347_), .A3(new_n344_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n388_), .A2(new_n384_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT4), .B1(new_n427_), .B2(KEYINPUT92), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n427_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n425_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n421_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n424_), .A2(new_n425_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT4), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n424_), .A2(new_n422_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n431_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n433_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n420_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n434_), .A2(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n369_), .A2(new_n414_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n331_), .A2(KEYINPUT96), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n322_), .A2(new_n323_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT98), .A4(new_n319_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n333_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n413_), .A2(new_n441_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n443_), .A2(new_n444_), .A3(new_n319_), .A4(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT97), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n318_), .A2(KEYINPUT27), .A3(new_n314_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(KEYINPUT96), .A2(new_n331_), .B1(new_n450_), .B2(new_n296_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n444_), .A4(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n295_), .A2(KEYINPUT32), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n328_), .A2(new_n300_), .A3(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n441_), .B(new_n455_), .C1(new_n289_), .C2(new_n454_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT93), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n432_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n420_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n429_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(KEYINPUT93), .A3(new_n420_), .A4(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT33), .B(new_n421_), .C1(new_n430_), .C2(new_n433_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n434_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n321_), .A2(new_n314_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n456_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n413_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n449_), .A2(new_n453_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n446_), .B1(new_n369_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n474_));
  OR2_X1    g273(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n419_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n474_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n482_), .A3(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n480_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n486_), .A3(new_n487_), .A4(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  XOR2_X1   g296(.A(G85gat), .B(G92gat), .Z(new_n498_));
  AND3_X1   g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n490_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G64gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G57gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n417_), .A2(G64gat), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT65), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT65), .B1(new_n503_), .B2(new_n504_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT11), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G71gat), .B(G78gat), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n417_), .A2(G64gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n502_), .A2(G57gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT11), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT65), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n509_), .B1(new_n507_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n501_), .B1(new_n511_), .B2(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n505_), .A2(new_n506_), .A3(KEYINPUT11), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n516_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n508_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n496_), .A2(new_n498_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n523_), .A2(new_n527_), .A3(new_n510_), .A4(new_n490_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n520_), .A2(new_n528_), .A3(KEYINPUT12), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n510_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n501_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n520_), .B2(new_n528_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G120gat), .B(G148gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT66), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT5), .B(G176gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n534_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n542_), .B1(new_n546_), .B2(new_n536_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n544_), .A2(KEYINPUT13), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT13), .B1(new_n544_), .B2(new_n547_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(G36gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(G29gat), .ZN(new_n554_));
  INV_X1    g353(.A(G29gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(G36gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT68), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G43gat), .B(G50gat), .Z(new_n560_));
  NOR3_X1   g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G43gat), .B(G50gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n554_), .A2(new_n556_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT68), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G1gat), .A2(G8gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT14), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(G1gat), .ZN(new_n572_));
  INV_X1    g371(.A(G8gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n569_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n571_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n567_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n571_), .B(new_n575_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n560_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n564_), .A2(new_n562_), .A3(new_n565_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n552_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n579_), .A2(new_n582_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT15), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n561_), .B2(new_n566_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT15), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n585_), .B1(new_n589_), .B2(new_n579_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n584_), .B1(new_n590_), .B2(new_n552_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G169gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n244_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n591_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n551_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n473_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n567_), .A2(new_n527_), .A3(new_n490_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT67), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT67), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(G232gat), .A3(G233gat), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT34), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n602_), .A2(new_n604_), .A3(KEYINPUT34), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT72), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT15), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT15), .B1(new_n580_), .B2(new_n581_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n501_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n607_), .A2(new_n615_), .A3(new_n608_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT69), .ZN(new_n617_));
  AND4_X1   g416(.A1(new_n600_), .A2(new_n611_), .A3(new_n614_), .A4(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT70), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n501_), .A2(new_n582_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT69), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n616_), .B(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n619_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n600_), .A2(KEYINPUT70), .A3(new_n617_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n614_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n610_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n618_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT71), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(G190gat), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(G218gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(G218gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT36), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n627_), .A2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n631_), .A2(KEYINPUT36), .A3(new_n632_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n633_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n627_), .B2(KEYINPUT73), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT73), .ZN(new_n638_));
  AOI211_X1 g437(.A(new_n638_), .B(new_n618_), .C1(new_n626_), .C2(new_n625_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n634_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n635_), .A2(new_n633_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n634_), .B(KEYINPUT37), .C1(new_n627_), .C2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G127gat), .B(G155gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT16), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(G183gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(new_n248_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT17), .ZN(new_n651_));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n579_), .B(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(new_n530_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT17), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n656_), .B2(new_n650_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n646_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT74), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n599_), .A2(new_n572_), .A3(new_n660_), .A4(new_n441_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT38), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n472_), .A2(new_n369_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n446_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n658_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n598_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n640_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n441_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n661_), .A2(new_n662_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n663_), .A2(new_n671_), .A3(new_n672_), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n599_), .A2(new_n660_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n333_), .A2(new_n445_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n674_), .A2(G8gat), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G8gat), .B1(new_n669_), .B2(new_n676_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n682_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n684_), .B(new_n677_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1325gat));
  OAI21_X1  g485(.A(G15gat), .B1(new_n669_), .B2(new_n369_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT41), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n674_), .A2(G15gat), .A3(new_n369_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1326gat));
  OAI21_X1  g489(.A(G22gat), .B1(new_n669_), .B2(new_n413_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n413_), .A2(G22gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n674_), .B2(new_n694_), .ZN(G1327gat));
  NOR2_X1   g494(.A1(new_n598_), .A2(new_n658_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n646_), .B2(KEYINPUT101), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n699_), .B1(new_n473_), .B2(new_n646_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n367_), .A2(new_n368_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n365_), .A2(new_n352_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n448_), .A2(KEYINPUT97), .B1(new_n470_), .B2(new_n413_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n453_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n645_), .B(new_n698_), .C1(new_n705_), .C2(new_n446_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n697_), .B1(new_n700_), .B2(new_n706_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n555_), .B(new_n670_), .C1(new_n707_), .C2(KEYINPUT44), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n707_), .A2(KEYINPUT44), .ZN(new_n709_));
  INV_X1    g508(.A(new_n640_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n667_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT102), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n597_), .B(new_n712_), .C1(new_n705_), .C2(new_n446_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT103), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n666_), .A2(new_n715_), .A3(new_n597_), .A4(new_n712_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(new_n716_), .A3(new_n441_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n708_), .A2(new_n709_), .B1(new_n555_), .B2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n676_), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n553_), .B1(new_n709_), .B2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n714_), .A2(new_n716_), .A3(new_n553_), .A4(new_n675_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n721_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n700_), .A2(new_n706_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n675_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n707_), .A2(KEYINPUT44), .ZN(new_n729_));
  OAI21_X1  g528(.A(G36gat), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n722_), .B(KEYINPUT45), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT46), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n725_), .A2(new_n732_), .ZN(G1329gat));
  NAND3_X1  g532(.A1(new_n714_), .A2(new_n716_), .A3(new_n703_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT104), .B(G43gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n727_), .A2(G43gat), .A3(new_n703_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n729_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT47), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(new_n736_), .C1(new_n737_), .C2(new_n729_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1330gat));
  INV_X1    g541(.A(G50gat), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n714_), .A2(new_n716_), .A3(new_n743_), .A4(new_n414_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n413_), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n709_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n747_), .B2(G50gat), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT105), .B(new_n743_), .C1(new_n709_), .C2(new_n746_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n744_), .B1(new_n748_), .B2(new_n749_), .ZN(G1331gat));
  NOR2_X1   g549(.A1(new_n473_), .A2(new_n710_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n550_), .A2(new_n595_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n667_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT106), .B1(new_n670_), .B2(new_n417_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(KEYINPUT106), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n757_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n666_), .A2(new_n660_), .A3(new_n752_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n441_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n758_), .B1(new_n762_), .B2(new_n417_), .ZN(G1332gat));
  OAI21_X1  g562(.A(G64gat), .B1(new_n755_), .B2(new_n676_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT48), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n502_), .A3(new_n675_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n755_), .B2(new_n369_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT49), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n369_), .A2(G71gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n760_), .B2(new_n770_), .ZN(G1334gat));
  OAI21_X1  g570(.A(G78gat), .B1(new_n755_), .B2(new_n413_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT50), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n413_), .A2(G78gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n760_), .B2(new_n774_), .ZN(G1335gat));
  OAI211_X1 g574(.A(new_n712_), .B(new_n752_), .C1(new_n705_), .C2(new_n446_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT107), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n666_), .A2(new_n778_), .A3(new_n712_), .A4(new_n752_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n419_), .A3(new_n441_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n726_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n753_), .A2(new_n658_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n782_), .A2(new_n670_), .A3(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n785_), .B2(new_n419_), .ZN(G1336gat));
  AOI21_X1  g585(.A(G92gat), .B1(new_n780_), .B2(new_n675_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n782_), .A2(new_n784_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n676_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(G1337gat));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n726_), .A2(new_n703_), .A3(new_n783_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G99gat), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n369_), .A2(new_n482_), .A3(new_n481_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n780_), .A2(KEYINPUT108), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT108), .B1(new_n780_), .B2(new_n794_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT51), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n793_), .B(new_n799_), .C1(new_n796_), .C2(new_n795_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1338gat));
  XNOR2_X1  g600(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n413_), .B(new_n784_), .C1(new_n700_), .C2(new_n706_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n493_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n726_), .A2(new_n414_), .A3(new_n783_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n413_), .A2(G106gat), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n803_), .B1(new_n809_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n812_), .B(KEYINPUT110), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(new_n802_), .A3(new_n806_), .A4(new_n808_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1339gat));
  NAND4_X1  g617(.A1(new_n333_), .A2(new_n703_), .A3(new_n441_), .A4(new_n445_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n595_), .A2(new_n544_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n529_), .A2(new_n545_), .A3(new_n532_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n824_));
  AOI211_X1 g623(.A(KEYINPUT55), .B(new_n545_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n822_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT113), .B1(new_n826_), .B2(new_n542_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n821_), .B1(new_n827_), .B2(KEYINPUT56), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829_));
  INV_X1    g628(.A(new_n822_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n535_), .A2(KEYINPUT55), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n546_), .A2(new_n823_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n833_), .B2(new_n543_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n828_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n577_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n585_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n579_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(KEYINPUT114), .A3(new_n578_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n552_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n578_), .A2(new_n583_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n594_), .B1(new_n845_), .B2(new_n552_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n591_), .A2(new_n594_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n547_), .B2(new_n544_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n710_), .B1(new_n837_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(KEYINPUT57), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n543_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n546_), .A2(new_n536_), .A3(new_n542_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT116), .B1(new_n849_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n544_), .A2(new_n859_), .A3(new_n848_), .A4(new_n847_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n826_), .A2(new_n835_), .A3(new_n542_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n856_), .A2(new_n861_), .A3(KEYINPUT58), .A4(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n856_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n864_), .A2(new_n865_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n852_), .A2(new_n855_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n850_), .B1(new_n828_), .B2(new_n836_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n854_), .B1(new_n868_), .B2(new_n710_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n658_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n548_), .A2(new_n549_), .A3(new_n595_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n642_), .A2(new_n871_), .A3(new_n658_), .A4(new_n644_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n872_), .B(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n413_), .B(new_n820_), .C1(new_n870_), .C2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n341_), .A3(new_n595_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n829_), .B(KEYINPUT56), .C1(new_n833_), .C2(new_n543_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n821_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n827_), .A2(KEYINPUT56), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n851_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n640_), .A3(new_n855_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n864_), .A2(new_n865_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n645_), .A3(new_n863_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n869_), .A2(new_n886_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n667_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n875_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n414_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n880_), .B1(new_n892_), .B2(new_n820_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n875_), .B1(new_n889_), .B2(new_n667_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n894_), .A2(KEYINPUT59), .A3(new_n414_), .A4(new_n819_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n879_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n876_), .A2(KEYINPUT59), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n892_), .A2(new_n880_), .A3(new_n820_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(KEYINPUT117), .A3(new_n898_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n896_), .A2(new_n899_), .A3(new_n595_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n878_), .B1(new_n900_), .B2(new_n341_), .ZN(G1340gat));
  NOR2_X1   g700(.A1(new_n550_), .A2(G120gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n877_), .B1(KEYINPUT60), .B2(new_n902_), .ZN(new_n903_));
  AND4_X1   g702(.A1(new_n551_), .A2(new_n903_), .A3(new_n897_), .A4(new_n898_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n904_), .A2(new_n334_), .B1(KEYINPUT60), .B2(new_n903_), .ZN(G1341gat));
  NAND3_X1  g704(.A1(new_n896_), .A2(new_n899_), .A3(new_n658_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(G127gat), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n667_), .A2(G127gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n876_), .B2(new_n908_), .ZN(G1342gat));
  NAND3_X1  g708(.A1(new_n896_), .A2(new_n899_), .A3(new_n645_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G134gat), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n876_), .A2(G134gat), .A3(new_n640_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n911_), .A2(KEYINPUT118), .A3(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1343gat));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n703_), .A2(new_n413_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n675_), .A2(new_n920_), .A3(new_n670_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n921_), .A2(KEYINPUT119), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(KEYINPUT119), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n918_), .B1(new_n924_), .B2(new_n894_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n894_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n922_), .A2(KEYINPUT120), .A3(new_n926_), .A4(new_n923_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n595_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n551_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT121), .B(G148gat), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n931_), .B(new_n932_), .Z(G1345gat));
  NAND2_X1  g732(.A1(new_n928_), .A2(new_n658_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT61), .B(G155gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1346gat));
  AOI21_X1  g735(.A(new_n640_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938_));
  OR3_X1    g737(.A1(new_n937_), .A2(new_n938_), .A3(G162gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n937_), .B2(G162gat), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n645_), .A2(G162gat), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n939_), .A2(new_n940_), .B1(new_n928_), .B2(new_n941_), .ZN(G1347gat));
  INV_X1    g741(.A(new_n892_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n675_), .A2(new_n703_), .A3(new_n670_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n595_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n236_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n946_), .A2(G169gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n947_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(new_n948_), .B2(new_n949_), .ZN(G1348gat));
  NAND2_X1  g750(.A1(new_n945_), .A2(new_n551_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G176gat), .ZN(G1349gat));
  OR4_X1    g752(.A1(new_n667_), .A2(new_n943_), .A3(new_n215_), .A4(new_n944_), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n954_), .A2(KEYINPUT124), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(KEYINPUT124), .ZN(new_n956_));
  AOI21_X1  g755(.A(G183gat), .B1(new_n945_), .B2(new_n658_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n945_), .A2(new_n710_), .A3(new_n272_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n943_), .A2(new_n646_), .A3(new_n944_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n960_), .B2(new_n212_), .ZN(G1351gat));
  NOR4_X1   g760(.A1(new_n894_), .A2(new_n441_), .A3(new_n676_), .A4(new_n920_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n962_), .A2(G197gat), .A3(new_n595_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n964_), .ZN(new_n966_));
  AOI21_X1  g765(.A(G197gat), .B1(new_n962_), .B2(new_n595_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n965_), .A2(new_n966_), .A3(new_n967_), .ZN(G1352gat));
  AND2_X1   g767(.A1(new_n962_), .A2(new_n551_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(new_n253_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n243_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n970_), .B1(KEYINPUT126), .B2(new_n971_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n972_), .B1(KEYINPUT126), .B2(new_n971_), .ZN(G1353gat));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n658_), .B1(new_n974_), .B2(new_n248_), .ZN(new_n975_));
  XOR2_X1   g774(.A(new_n975_), .B(KEYINPUT127), .Z(new_n976_));
  NAND2_X1  g775(.A1(new_n962_), .A2(new_n976_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n974_), .A2(new_n248_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n977_), .B(new_n978_), .ZN(G1354gat));
  NAND3_X1  g778(.A1(new_n962_), .A2(new_n246_), .A3(new_n710_), .ZN(new_n980_));
  AND2_X1   g779(.A1(new_n962_), .A2(new_n645_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n980_), .B1(new_n981_), .B2(new_n246_), .ZN(G1355gat));
endmodule


