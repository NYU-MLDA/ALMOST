//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT30), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT24), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT78), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n206_), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n207_), .A2(new_n208_), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n216_), .A2(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT22), .B1(new_n207_), .B2(KEYINPUT79), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n208_), .B(new_n225_), .C1(new_n226_), .C2(KEYINPUT79), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n212_), .B(new_n213_), .C1(G183gat), .C2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G71gat), .B(G99gat), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n232_), .B(G43gat), .Z(new_n233_));
  NOR2_X1   g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n233_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n205_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n205_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n238_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT81), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G134gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G127gat), .ZN(new_n251_));
  INV_X1    g050(.A(G127gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G134gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n251_), .A2(new_n253_), .A3(new_n248_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n246_), .B1(new_n249_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT80), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n247_), .A2(new_n248_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(new_n245_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT31), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n242_), .A2(new_n244_), .A3(new_n261_), .ZN(new_n262_));
  OR4_X1    g061(.A1(new_n243_), .A2(new_n240_), .A3(new_n237_), .A4(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT1), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT82), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(KEYINPUT82), .B(new_n267_), .C1(new_n268_), .C2(KEYINPUT1), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n267_), .A2(KEYINPUT1), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(KEYINPUT3), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n275_), .B(KEYINPUT2), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n267_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(new_n268_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n274_), .A2(new_n278_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT90), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n255_), .A2(new_n286_), .A3(new_n259_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n284_), .B(new_n285_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n274_), .A2(new_n278_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n281_), .A2(new_n283_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n260_), .A2(KEYINPUT90), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n255_), .A2(new_n286_), .A3(new_n259_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n255_), .A2(new_n259_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT91), .B1(new_n296_), .B2(new_n284_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n266_), .B(new_n289_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n299_), .A3(new_n260_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n289_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(KEYINPUT4), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n298_), .B1(new_n303_), .B2(new_n266_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G85gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT0), .B(G57gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n310_), .B(new_n298_), .C1(new_n303_), .C2(new_n266_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(G197gat), .A2(G204gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G197gat), .A2(G204gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(KEYINPUT21), .A3(new_n314_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G211gat), .B(G218gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G169gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT88), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n208_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n229_), .B(KEYINPUT87), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n228_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n322_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n220_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n214_), .B1(new_n220_), .B2(new_n331_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n330_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n216_), .A2(new_n217_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n218_), .A2(new_n219_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT85), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n338_), .A2(KEYINPUT86), .A3(new_n332_), .A4(new_n214_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n329_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT19), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n231_), .A2(new_n322_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n340_), .A2(KEYINPUT20), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G8gat), .B(G36gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n231_), .B2(new_n322_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n325_), .A2(new_n328_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n335_), .A2(new_n352_), .A3(new_n339_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n353_), .B2(new_n322_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n345_), .B(new_n350_), .C1(new_n354_), .C2(new_n343_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n323_), .A2(KEYINPUT88), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n323_), .A2(KEYINPUT88), .ZN(new_n358_));
  AOI21_X1  g157(.A(G176gat), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n320_), .B(new_n321_), .C1(new_n359_), .C2(new_n327_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n333_), .A2(new_n334_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n344_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n338_), .A2(new_n332_), .A3(new_n214_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n329_), .B2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(KEYINPUT93), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n342_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n354_), .A2(new_n343_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n350_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n356_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n312_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT94), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n309_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n345_), .B1(new_n354_), .B2(new_n343_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n349_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n345_), .B(new_n349_), .C1(new_n354_), .C2(new_n343_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(KEYINPUT89), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n378_), .A2(new_n383_), .A3(new_n379_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n303_), .A2(new_n266_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n303_), .A2(KEYINPUT92), .A3(new_n266_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n266_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n308_), .B1(new_n302_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n304_), .A2(KEYINPUT33), .A3(new_n308_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n377_), .A2(new_n385_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n312_), .A2(new_n395_), .A3(new_n373_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n375_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n322_), .B1(new_n284_), .B2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G22gat), .B(G50gat), .Z(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n403_));
  NOR3_X1   g202(.A1(new_n292_), .A2(KEYINPUT29), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n284_), .B2(new_n398_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT84), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n412_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n402_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n413_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n401_), .A3(new_n414_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n397_), .A2(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n367_), .A2(KEYINPUT93), .B1(new_n322_), .B2(new_n231_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n362_), .A2(new_n363_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n343_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n354_), .A2(new_n343_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n379_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n354_), .A2(new_n343_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT95), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n349_), .A4(new_n345_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n381_), .A2(KEYINPUT95), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n425_), .A2(new_n428_), .A3(KEYINPUT27), .A4(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT96), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n371_), .B2(new_n379_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(KEYINPUT96), .A3(new_n429_), .A4(new_n428_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n385_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n432_), .A2(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n312_), .A2(new_n419_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n265_), .B1(new_n420_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT98), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n432_), .A2(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n437_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n419_), .A2(new_n263_), .A3(new_n262_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(new_n312_), .ZN(new_n446_));
  AND4_X1   g245(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .A4(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n442_), .B1(new_n438_), .B2(new_n446_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n441_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G8gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT76), .ZN(new_n452_));
  INV_X1    g251(.A(G22gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n203_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G15gat), .A2(G22gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G1gat), .A2(G8gat), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n454_), .A2(new_n455_), .B1(KEYINPUT14), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n452_), .B(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G29gat), .B(G36gat), .Z(new_n459_));
  XOR2_X1   g258(.A(G43gat), .B(G50gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n461_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT77), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OR3_X1    g265(.A1(new_n458_), .A2(KEYINPUT77), .A3(new_n461_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n458_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n461_), .B(KEYINPUT15), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n465_), .A3(new_n463_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G113gat), .B(G141gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(G169gat), .B(G197gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n450_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT10), .B(G99gat), .Z(new_n479_));
  INV_X1    g278(.A(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G99gat), .A3(G106gat), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n479_), .A2(new_n480_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(G85gat), .A2(G92gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(KEYINPUT9), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT9), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT66), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT9), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n487_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n488_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  AOI211_X1 g294(.A(KEYINPUT67), .B(new_n487_), .C1(new_n490_), .C2(new_n492_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n485_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n482_), .A2(new_n484_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n500_));
  INV_X1    g299(.A(G99gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n480_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT8), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n487_), .A2(new_n486_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n497_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT69), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n512_), .B2(KEYINPUT11), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n515_));
  XOR2_X1   g314(.A(G71gat), .B(G78gat), .Z(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n511_), .A3(KEYINPUT11), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(KEYINPUT11), .B2(new_n512_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n517_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n513_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n497_), .B(KEYINPUT68), .C1(new_n506_), .C2(new_n507_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n510_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n508_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n482_), .A2(new_n484_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n502_), .A2(new_n499_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n505_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT8), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(KEYINPUT70), .A3(new_n497_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n518_), .A2(KEYINPUT12), .A3(new_n521_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n524_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G230gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n522_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n523_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT68), .B1(new_n532_), .B2(new_n497_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n536_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n524_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n539_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT5), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n546_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n557_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(KEYINPUT13), .A3(new_n555_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n526_), .A2(new_n470_), .A3(new_n533_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n510_), .A2(new_n461_), .A3(new_n523_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n566_), .A2(new_n567_), .A3(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(new_n571_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n566_), .A2(new_n567_), .A3(new_n576_), .A4(new_n572_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT36), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT73), .Z(new_n586_));
  NAND3_X1  g385(.A1(new_n575_), .A2(new_n577_), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n565_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n582_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT74), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n578_), .B2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n575_), .A2(KEYINPUT74), .A3(new_n577_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n588_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n522_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n458_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n604_), .A2(new_n605_), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n600_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n597_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n564_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n478_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT99), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n478_), .A2(new_n616_), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(KEYINPUT100), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  INV_X1    g422(.A(new_n312_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(G1gat), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n622_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n450_), .A2(new_n594_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n477_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n563_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n610_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n624_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n623_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n633_), .A3(new_n634_), .ZN(G1324gat));
  NOR2_X1   g434(.A1(new_n438_), .A2(G8gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n620_), .A2(new_n621_), .A3(new_n636_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n397_), .A2(new_n419_), .B1(new_n439_), .B2(new_n438_), .ZN(new_n638_));
  OAI22_X1  g437(.A1(new_n638_), .A2(new_n265_), .B1(new_n448_), .B2(new_n447_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n438_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n594_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .A4(new_n630_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G8gat), .B1(new_n642_), .B2(new_n643_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT102), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n642_), .A2(new_n643_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(G8gat), .A4(new_n644_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n647_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n637_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  AOI21_X1  g455(.A(new_n203_), .B1(new_n631_), .B2(new_n265_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT41), .ZN(new_n658_));
  INV_X1    g457(.A(new_n618_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n203_), .A3(new_n265_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1326gat));
  INV_X1    g460(.A(new_n419_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n453_), .B1(new_n631_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT42), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n659_), .A2(new_n453_), .A3(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n594_), .A2(new_n610_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n564_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n478_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n312_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n629_), .A2(new_n611_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n597_), .B1(new_n639_), .B2(KEYINPUT103), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675_));
  OAI221_X1 g474(.A(new_n675_), .B1(new_n447_), .B2(new_n448_), .C1(new_n638_), .C2(new_n265_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n597_), .A2(KEYINPUT43), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n639_), .A2(KEYINPUT104), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n672_), .B1(new_n677_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n672_), .C1(new_n677_), .C2(new_n683_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n312_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n671_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n686_), .A2(new_n640_), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n438_), .B(KEYINPUT105), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n669_), .A2(G36gat), .A3(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n692_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n692_), .A2(KEYINPUT46), .A3(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1329gat));
  NAND4_X1  g500(.A1(new_n686_), .A2(G43gat), .A3(new_n265_), .A4(new_n687_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT107), .B(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n669_), .B2(new_n264_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g505(.A1(new_n669_), .A2(G50gat), .A3(new_n419_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n686_), .A2(new_n662_), .A3(new_n687_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT108), .ZN(new_n709_));
  OAI21_X1  g508(.A(G50gat), .B1(new_n708_), .B2(KEYINPUT108), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(G1331gat));
  NAND2_X1  g510(.A1(new_n639_), .A2(new_n477_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n712_), .A2(KEYINPUT109), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(KEYINPUT109), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n612_), .A2(new_n563_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n312_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n628_), .A2(new_n610_), .ZN(new_n722_));
  AND4_X1   g521(.A1(new_n639_), .A2(new_n564_), .A3(new_n641_), .A4(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n312_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n720_), .B2(new_n724_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n693_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n723_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n726_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n718_), .B2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n723_), .B2(new_n265_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT49), .Z(new_n735_));
  NAND4_X1  g534(.A1(new_n716_), .A2(new_n733_), .A3(new_n265_), .A4(new_n717_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT111), .Z(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n723_), .B2(new_n662_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT50), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n662_), .A2(new_n739_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n718_), .B2(new_n742_), .ZN(G1335gat));
  OR2_X1    g542(.A1(new_n563_), .A2(new_n667_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n715_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n312_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n563_), .A2(new_n628_), .A3(new_n611_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n677_), .B2(new_n683_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT103), .B1(new_n441_), .B2(new_n449_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n676_), .A3(new_n596_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT43), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n639_), .A2(KEYINPUT104), .A3(new_n678_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT104), .B1(new_n639_), .B2(new_n678_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n756_), .A3(KEYINPUT112), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n748_), .B1(new_n750_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n312_), .A2(G85gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT113), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n746_), .B1(new_n758_), .B2(new_n760_), .ZN(G1336gat));
  INV_X1    g560(.A(G92gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n745_), .A2(new_n762_), .A3(new_n640_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n758_), .A2(new_n727_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n762_), .ZN(G1337gat));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(KEYINPUT51), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(KEYINPUT51), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n501_), .B1(new_n758_), .B2(new_n265_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n265_), .A2(new_n479_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n715_), .A2(new_n744_), .A3(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n767_), .B(new_n768_), .C1(new_n769_), .C2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n677_), .A2(new_n683_), .A3(new_n749_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT112), .B1(new_n753_), .B2(new_n756_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n265_), .B(new_n747_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G99gat), .ZN(new_n776_));
  INV_X1    g575(.A(new_n771_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n776_), .A2(new_n766_), .A3(KEYINPUT51), .A4(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n772_), .A2(new_n778_), .ZN(G1338gat));
  NAND2_X1  g578(.A1(new_n662_), .A2(new_n480_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n715_), .A2(new_n744_), .A3(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n662_), .B(new_n747_), .C1(new_n677_), .C2(new_n683_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n782_), .B2(G106gat), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n747_), .A2(new_n662_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n753_), .B2(new_n756_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n788_), .B2(new_n480_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(KEYINPUT52), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n785_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n785_), .B2(new_n791_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796_));
  INV_X1    g595(.A(new_n473_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n465_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n476_), .B1(new_n471_), .B2(new_n799_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n797_), .A2(new_n476_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n558_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n522_), .B1(new_n510_), .B2(new_n523_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n524_), .B(new_n535_), .C1(new_n804_), .C2(KEYINPUT12), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n805_), .B2(new_n548_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n548_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n536_), .A2(new_n545_), .A3(KEYINPUT55), .A4(new_n539_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n553_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(new_n813_), .A3(new_n553_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n811_), .A2(KEYINPUT119), .A3(new_n812_), .A4(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n477_), .A2(new_n556_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n553_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n810_), .B2(KEYINPUT118), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n814_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n802_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n796_), .B1(new_n823_), .B2(new_n641_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n801_), .A2(new_n555_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n810_), .A2(new_n812_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n818_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n596_), .B1(new_n830_), .B2(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT121), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n596_), .C1(new_n830_), .C2(KEYINPUT58), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n610_), .B1(new_n827_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n563_), .A2(KEYINPUT117), .A3(new_n722_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n722_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n839_), .B1(new_n844_), .B2(new_n597_), .ZN(new_n845_));
  AOI211_X1 g644(.A(KEYINPUT54), .B(new_n596_), .C1(new_n840_), .C2(new_n843_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n838_), .A2(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n640_), .A2(new_n624_), .A3(new_n445_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT59), .ZN(new_n852_));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852_), .B2(new_n477_), .ZN(new_n853_));
  OR3_X1    g652(.A1(new_n851_), .A2(G113gat), .A3(new_n477_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n852_), .B2(new_n563_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT60), .ZN(new_n857_));
  AOI21_X1  g656(.A(G120gat), .B1(new_n564_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT122), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n857_), .B2(G120gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n859_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n856_), .B1(new_n851_), .B2(new_n862_), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n852_), .B2(new_n610_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n851_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n252_), .A3(new_n611_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1342gat));
  OAI21_X1  g666(.A(G134gat), .B1(new_n852_), .B2(new_n597_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n250_), .A3(new_n594_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1343gat));
  AOI21_X1  g669(.A(new_n265_), .B1(new_n838_), .B2(new_n848_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n693_), .A2(new_n662_), .A3(new_n312_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT123), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n811_), .A2(new_n812_), .A3(new_n814_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n815_), .B(new_n816_), .C1(new_n875_), .C2(new_n820_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n594_), .B1(new_n876_), .B2(new_n802_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT57), .B1(new_n877_), .B2(new_n796_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n826_), .A3(new_n836_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n847_), .B1(new_n879_), .B2(new_n610_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n880_), .A2(new_n881_), .A3(new_n265_), .A4(new_n872_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n628_), .B1(new_n874_), .B2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n835_), .A2(new_n833_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886_));
  INV_X1    g685(.A(new_n818_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n553_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n886_), .B1(new_n889_), .B2(new_n828_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n834_), .B1(new_n890_), .B2(new_n596_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n885_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n823_), .A2(new_n641_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT120), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n894_), .B2(KEYINPUT57), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n611_), .B1(new_n895_), .B2(new_n826_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n264_), .B(new_n873_), .C1(new_n896_), .C2(new_n847_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n881_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n871_), .A2(KEYINPUT123), .A3(new_n873_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n563_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT124), .B(G148gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1345gat));
  AOI21_X1  g701(.A(new_n610_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  INV_X1    g704(.A(G162gat), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n906_), .B(new_n597_), .C1(new_n898_), .C2(new_n899_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n641_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n908_), .B2(G162gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n594_), .B1(new_n874_), .B2(new_n882_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(new_n906_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n907_), .B1(new_n909_), .B2(new_n912_), .ZN(G1347gat));
  OAI211_X1 g712(.A(new_n446_), .B(new_n727_), .C1(new_n896_), .C2(new_n847_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n477_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT127), .B1(new_n915_), .B2(new_n207_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n917_), .B(G169gat), .C1(new_n914_), .C2(new_n477_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n919_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT127), .B(new_n921_), .C1(new_n915_), .C2(new_n207_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n915_), .A2(new_n324_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(new_n922_), .A3(new_n923_), .ZN(G1348gat));
  NOR2_X1   g723(.A1(new_n914_), .A2(new_n563_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n208_), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n914_), .A2(new_n610_), .ZN(new_n927_));
  MUX2_X1   g726(.A(G183gat), .B(new_n216_), .S(new_n927_), .Z(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n914_), .B2(new_n597_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n594_), .A2(new_n217_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n914_), .B2(new_n930_), .ZN(G1351gat));
  AND3_X1   g730(.A1(new_n871_), .A2(new_n439_), .A3(new_n727_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n628_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n564_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g735(.A(KEYINPUT63), .B(G211gat), .C1(new_n932_), .C2(new_n611_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n932_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n610_), .ZN(new_n939_));
  XOR2_X1   g738(.A(KEYINPUT63), .B(G211gat), .Z(new_n940_));
  AOI21_X1  g739(.A(new_n937_), .B1(new_n939_), .B2(new_n940_), .ZN(G1354gat));
  OR3_X1    g740(.A1(new_n938_), .A2(G218gat), .A3(new_n641_), .ZN(new_n942_));
  OAI21_X1  g741(.A(G218gat), .B1(new_n938_), .B2(new_n597_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1355gat));
endmodule


