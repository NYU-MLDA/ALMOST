//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT75), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT23), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n214_), .B1(KEYINPUT77), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(KEYINPUT77), .B2(new_n217_), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n204_), .B(KEYINPUT76), .C1(new_n207_), .C2(new_n208_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n211_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n213_), .A2(KEYINPUT79), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(KEYINPUT79), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n217_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n207_), .B1(KEYINPUT78), .B2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n228_), .B(new_n232_), .C1(KEYINPUT78), .C2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n222_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT31), .Z(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n222_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G71gat), .B(G99gat), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n241_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n243_), .A3(new_n239_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(KEYINPUT82), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n247_), .A2(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n250_), .B1(new_n253_), .B2(KEYINPUT82), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT83), .B1(new_n259_), .B2(new_n250_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n256_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n257_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n246_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n260_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n259_), .A2(new_n250_), .A3(KEYINPUT83), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT80), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n256_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n266_), .A2(G227gat), .A3(G233gat), .A4(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G15gat), .B(G43gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n263_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n245_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n263_), .A2(new_n268_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n269_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n242_), .A2(new_n244_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n263_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G197gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(G204gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT21), .B1(new_n283_), .B2(KEYINPUT88), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n281_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(KEYINPUT89), .ZN(new_n289_));
  INV_X1    g088(.A(new_n285_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT89), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n289_), .A2(KEYINPUT21), .A3(new_n290_), .A4(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT90), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT87), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n294_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT2), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(KEYINPUT86), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n299_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(KEYINPUT86), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n305_), .A2(new_n306_), .B1(new_n307_), .B2(KEYINPUT3), .ZN(new_n308_));
  OR4_X1    g107(.A1(new_n307_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n309_));
  INV_X1    g108(.A(G141gat), .ZN(new_n310_));
  INV_X1    g109(.A(G148gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n307_), .B2(KEYINPUT3), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n304_), .A2(new_n308_), .A3(new_n309_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  OR2_X1    g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n305_), .B1(new_n318_), .B2(new_n312_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n316_), .ZN(new_n322_));
  OAI221_X1 g121(.A(new_n319_), .B1(new_n318_), .B2(new_n312_), .C1(new_n320_), .C2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT29), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n298_), .A2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(G228gat), .B(G233gat), .C1(new_n295_), .C2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n325_), .A2(KEYINPUT87), .A3(new_n297_), .A4(new_n294_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G78gat), .B(G106gat), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(new_n330_), .A3(new_n328_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n324_), .A2(KEYINPUT29), .ZN(new_n335_));
  XOR2_X1   g134(.A(G22gat), .B(G50gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT28), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n330_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT91), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n332_), .A2(new_n340_), .A3(new_n333_), .A4(new_n338_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n279_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n345_));
  INV_X1    g144(.A(new_n294_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n222_), .A3(new_n233_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT20), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n351_));
  INV_X1    g150(.A(new_n208_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n202_), .A2(new_n203_), .B1(new_n352_), .B2(new_n205_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n225_), .A2(new_n220_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT93), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT93), .B1(new_n225_), .B2(new_n220_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT94), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT94), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n353_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n219_), .A2(new_n227_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n207_), .B1(new_n230_), .B2(new_n229_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n359_), .A2(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n350_), .B(new_n351_), .C1(new_n364_), .C2(new_n346_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n362_), .A2(new_n363_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n354_), .B(new_n355_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n360_), .B1(new_n370_), .B2(new_n353_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n361_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n346_), .B(new_n369_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT95), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT95), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n364_), .A2(new_n375_), .A3(new_n346_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n234_), .A2(new_n294_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n367_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n377_), .A2(KEYINPUT20), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  INV_X1    g180(.A(G92gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT18), .B(G64gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n368_), .A2(new_n380_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n368_), .B2(new_n380_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n345_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n317_), .A2(new_n323_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n324_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(KEYINPUT96), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT4), .B1(new_n391_), .B2(new_n392_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n324_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n395_), .B1(new_n401_), .B2(KEYINPUT97), .ZN(new_n402_));
  INV_X1    g201(.A(new_n396_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n390_), .A2(new_n253_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n391_), .A2(KEYINPUT4), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n403_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT97), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410_));
  INV_X1    g209(.A(G85gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G57gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  NOR3_X1   g213(.A1(new_n402_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n414_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n393_), .A2(new_n394_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n401_), .A2(KEYINPUT97), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n369_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n294_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n423_), .A2(new_n378_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n295_), .A2(new_n369_), .A3(new_n358_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT20), .A3(new_n377_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n367_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n385_), .B(KEYINPUT98), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n368_), .A2(new_n380_), .A3(new_n386_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(KEYINPUT27), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n344_), .A2(new_n389_), .A3(new_n421_), .A4(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT100), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n389_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n342_), .A2(new_n343_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n386_), .A2(KEYINPUT32), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n368_), .A2(new_n380_), .A3(new_n438_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n440_), .B(new_n441_), .C1(new_n415_), .C2(new_n420_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n436_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n418_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n418_), .A2(KEYINPUT33), .A3(new_n416_), .A4(new_n419_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n394_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n416_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n388_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n431_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n442_), .B(new_n443_), .C1(new_n451_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n279_), .ZN(new_n455_));
  AND4_X1   g254(.A1(KEYINPUT99), .A2(new_n437_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n414_), .B1(new_n402_), .B2(new_n409_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n439_), .B1(new_n457_), .B2(new_n444_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n436_), .B1(new_n458_), .B2(new_n441_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n387_), .A2(new_n388_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n460_), .A2(new_n447_), .A3(new_n450_), .A4(new_n446_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n279_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT99), .B1(new_n462_), .B2(new_n437_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n434_), .B1(new_n456_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT65), .ZN(new_n465_));
  AND2_X1   g264(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n466_));
  NOR2_X1   g265(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(G99gat), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n470_), .A2(KEYINPUT10), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(KEYINPUT10), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n479_), .A2(KEYINPUT9), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n411_), .A2(new_n382_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT9), .A3(new_n479_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n473_), .A2(new_n478_), .A3(new_n480_), .A4(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT7), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n470_), .A3(new_n469_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n476_), .A3(new_n477_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT8), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n481_), .A2(new_n479_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n483_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G57gat), .ZN(new_n493_));
  INV_X1    g292(.A(G64gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G57gat), .A2(G64gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G78gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT11), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n495_), .A2(new_n501_), .A3(new_n496_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n468_), .B1(new_n492_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n467_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n492_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n487_), .A2(new_n489_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT8), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n483_), .A3(new_n505_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n492_), .A2(new_n506_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT64), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n473_), .A2(new_n480_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n478_), .A2(new_n482_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n513_), .A2(new_n514_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(KEYINPUT64), .A3(new_n505_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n509_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n465_), .B1(new_n517_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n465_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n529_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n529_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(new_n527_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT13), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(KEYINPUT13), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G1gat), .B(G8gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT73), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547_));
  INV_X1    g346(.A(G1gat), .ZN(new_n548_));
  INV_X1    g347(.A(G8gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT14), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n546_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n546_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT68), .B(G43gat), .ZN(new_n555_));
  INV_X1    g354(.A(G50gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G29gat), .A2(G36gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(G29gat), .A2(G36gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n556_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(G29gat), .ZN(new_n561_));
  INV_X1    g360(.A(G36gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(G50gat), .A3(new_n557_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n555_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n564_), .A3(new_n555_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n554_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n573_));
  INV_X1    g372(.A(new_n567_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n565_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(KEYINPUT15), .A3(new_n567_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n554_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n554_), .A2(new_n568_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n570_), .A3(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G169gat), .B(G197gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n581_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n544_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n464_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n515_), .A2(new_n568_), .A3(new_n483_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n577_), .B2(new_n523_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT34), .Z(new_n593_));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n597_), .B2(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n590_), .A2(KEYINPUT69), .A3(new_n596_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT69), .B1(new_n590_), .B2(new_n596_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n600_), .B(new_n605_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT71), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n600_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n603_), .B(KEYINPUT36), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n610_), .A2(KEYINPUT37), .A3(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n608_), .A2(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(KEYINPUT72), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT72), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n618_), .A3(new_n612_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n619_), .A3(new_n608_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n621_), .B2(KEYINPUT37), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT74), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n554_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(new_n505_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628_));
  INV_X1    g427(.A(G211gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT16), .B(G183gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(KEYINPUT17), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT17), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n627_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n627_), .A2(new_n633_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n622_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n588_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n421_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n548_), .A3(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n620_), .B(KEYINPUT102), .Z(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n637_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n588_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(new_n640_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n643_), .B(new_n644_), .C1(new_n548_), .C2(new_n649_), .ZN(G1324gat));
  XNOR2_X1  g449(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n389_), .A2(new_n432_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n464_), .A2(new_n587_), .A3(new_n653_), .A4(new_n647_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(G8gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(KEYINPUT103), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n652_), .A3(G8gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(KEYINPUT103), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n639_), .A2(new_n549_), .A3(new_n653_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n651_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n658_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n661_), .B(new_n651_), .C1(new_n663_), .C2(new_n656_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1325gat));
  NAND2_X1  g465(.A1(new_n648_), .A2(new_n279_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G15gat), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT41), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT41), .ZN(new_n670_));
  INV_X1    g469(.A(G15gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n639_), .A2(new_n671_), .A3(new_n279_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n648_), .B2(new_n436_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT42), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n639_), .A2(new_n674_), .A3(new_n436_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(new_n637_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n620_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n588_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n561_), .A3(new_n640_), .ZN(new_n683_));
  OR2_X1    g482(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n684_));
  NAND2_X1  g483(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n433_), .B(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n437_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n462_), .A2(KEYINPUT99), .A3(new_n437_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT37), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n693_), .A2(new_n620_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n684_), .B(new_n685_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n464_), .A2(KEYINPUT105), .A3(KEYINPUT43), .A4(new_n622_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n544_), .A2(new_n586_), .A3(new_n679_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n695_), .A2(new_n696_), .A3(KEYINPUT44), .A4(new_n697_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(new_n640_), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n683_), .B1(new_n702_), .B2(new_n561_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n700_), .A2(new_n653_), .A3(new_n701_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n653_), .A2(KEYINPUT106), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n653_), .A2(KEYINPUT106), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(G36gat), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n464_), .A2(new_n587_), .A3(new_n680_), .A4(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(KEYINPUT45), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(KEYINPUT45), .ZN(new_n716_));
  OAI22_X1  g515(.A1(new_n715_), .A2(new_n716_), .B1(KEYINPUT107), .B2(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n707_), .B1(new_n709_), .B2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n706_), .B(new_n717_), .C1(new_n708_), .C2(G36gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n700_), .A2(new_n279_), .A3(new_n701_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G43gat), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n681_), .A2(G43gat), .A3(new_n455_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n722_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n722_), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n725_), .B(new_n728_), .C1(new_n723_), .C2(G43gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1330gat));
  NAND3_X1  g529(.A1(new_n682_), .A2(new_n556_), .A3(new_n436_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n700_), .A2(new_n436_), .A3(new_n701_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n556_), .ZN(G1331gat));
  NAND2_X1  g532(.A1(new_n544_), .A2(new_n586_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n692_), .A2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n638_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n640_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n735_), .A2(new_n647_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n421_), .A2(new_n493_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(G1332gat));
  INV_X1    g539(.A(new_n712_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n494_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT48), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n736_), .A2(new_n494_), .A3(new_n741_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n736_), .A2(new_n746_), .A3(new_n279_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n738_), .B2(new_n279_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n749_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n738_), .B2(new_n436_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT50), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n736_), .A2(new_n753_), .A3(new_n436_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1335gat));
  AND2_X1   g556(.A1(new_n735_), .A2(new_n680_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n640_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n734_), .A2(new_n679_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n695_), .A2(new_n696_), .A3(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n421_), .A2(new_n411_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  AOI21_X1  g562(.A(G92gat), .B1(new_n758_), .B2(new_n653_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n712_), .A2(new_n382_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  NAND4_X1  g565(.A1(new_n695_), .A2(new_n696_), .A3(new_n279_), .A4(new_n760_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n471_), .A2(new_n472_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n455_), .A2(new_n768_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n767_), .A2(G99gat), .B1(new_n758_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(KEYINPUT51), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n771_), .A2(KEYINPUT51), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n758_), .A2(new_n469_), .A3(new_n436_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n695_), .A2(new_n696_), .A3(new_n436_), .A4(new_n760_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n776_), .B(new_n782_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n511_), .A2(new_n516_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n525_), .B1(new_n787_), .B2(new_n507_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT113), .ZN(new_n790_));
  INV_X1    g589(.A(new_n517_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(new_n792_), .A3(KEYINPUT55), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n505_), .B1(new_n515_), .B2(new_n483_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n511_), .B(new_n516_), .C1(new_n796_), .C2(new_n468_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT113), .B(new_n795_), .C1(new_n797_), .C2(new_n525_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n792_), .B1(new_n788_), .B2(KEYINPUT55), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n517_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n794_), .A2(new_n800_), .A3(new_n536_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT56), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n794_), .A2(new_n800_), .A3(new_n803_), .A4(new_n536_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n802_), .A2(new_n535_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n578_), .A2(new_n571_), .A3(new_n579_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n584_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n581_), .A2(new_n584_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n805_), .A2(KEYINPUT116), .A3(KEYINPUT58), .A4(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n802_), .A2(new_n535_), .A3(new_n804_), .A4(new_n808_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n694_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n809_), .B(new_n813_), .C1(new_n814_), .C2(KEYINPUT115), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n816_), .B(new_n694_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n539_), .A2(new_n819_), .A3(new_n808_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n539_), .B2(new_n808_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n535_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n801_), .B2(KEYINPUT56), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n585_), .A3(new_n804_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n818_), .B1(new_n826_), .B2(new_n620_), .ZN(new_n827_));
  AOI211_X1 g626(.A(KEYINPUT57), .B(new_n621_), .C1(new_n822_), .C2(new_n825_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n815_), .A2(new_n817_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(new_n637_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n638_), .A2(new_n543_), .A3(new_n586_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n344_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n653_), .A2(new_n836_), .A3(new_n421_), .ZN(new_n837_));
  XOR2_X1   g636(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n585_), .A2(G113gat), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n829_), .A2(new_n841_), .ZN(new_n842_));
  OAI221_X1 g641(.A(KEYINPUT117), .B1(new_n827_), .B2(new_n828_), .C1(new_n815_), .C2(new_n817_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n637_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n833_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n845_), .A2(new_n837_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n839_), .B(new_n840_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n846_), .B2(new_n585_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1340gat));
  OAI21_X1  g650(.A(new_n839_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852_), .B2(new_n543_), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n543_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n846_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1341gat));
  AND2_X1   g656(.A1(new_n679_), .A2(G127gat), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n839_), .B(new_n858_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G127gat), .B1(new_n846_), .B2(new_n679_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  AND2_X1   g661(.A1(new_n622_), .A2(G134gat), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n839_), .B(new_n863_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G134gat), .B1(new_n846_), .B2(new_n646_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n443_), .A2(new_n421_), .A3(new_n279_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n712_), .A2(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT119), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n845_), .A2(KEYINPUT120), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n679_), .B1(new_n829_), .B2(new_n841_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n834_), .B1(new_n873_), .B2(new_n843_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n870_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n871_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n585_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n544_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n679_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  AOI21_X1  g683(.A(G162gat), .B1(new_n877_), .B2(new_n646_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n622_), .A2(G162gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT121), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n871_), .B2(new_n876_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT122), .B1(new_n885_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n877_), .A2(new_n887_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n645_), .B1(new_n871_), .B2(new_n876_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n892_), .C1(G162gat), .C2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n890_), .A2(new_n894_), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n830_), .A2(new_n834_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n712_), .A2(new_n640_), .A3(new_n836_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n896_), .A2(KEYINPUT124), .A3(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT124), .B1(new_n896_), .B2(new_n898_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n585_), .A3(new_n229_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n585_), .B(new_n897_), .C1(new_n830_), .C2(new_n834_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G169gat), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n906_), .A3(KEYINPUT62), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(KEYINPUT62), .B2(new_n905_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n905_), .B2(KEYINPUT62), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n903_), .B1(new_n908_), .B2(new_n909_), .ZN(G1348gat));
  NOR4_X1   g709(.A1(new_n874_), .A2(new_n230_), .A3(new_n543_), .A4(new_n898_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n902_), .A2(new_n544_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n230_), .ZN(G1349gat));
  NOR3_X1   g712(.A1(new_n901_), .A2(new_n202_), .A3(new_n637_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n835_), .A2(new_n679_), .A3(new_n897_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n915_), .A2(KEYINPUT125), .ZN(new_n916_));
  AOI21_X1  g715(.A(G183gat), .B1(new_n915_), .B2(KEYINPUT125), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n914_), .B1(new_n916_), .B2(new_n917_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n901_), .B2(new_n694_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n646_), .A2(new_n203_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n901_), .B2(new_n920_), .ZN(G1351gat));
  NOR4_X1   g720(.A1(new_n712_), .A2(new_n443_), .A3(new_n640_), .A4(new_n279_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n845_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n586_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n282_), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n543_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1353gat));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n845_), .A2(new_n922_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n637_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n932_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT127), .B1(new_n923_), .B2(new_n934_), .ZN(new_n935_));
  AND4_X1   g734(.A1(new_n929_), .A2(new_n933_), .A3(new_n629_), .A4(new_n935_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n933_), .A2(new_n935_), .B1(new_n929_), .B2(new_n629_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1354gat));
  AND3_X1   g737(.A1(new_n930_), .A2(G218gat), .A3(new_n622_), .ZN(new_n939_));
  AOI21_X1  g738(.A(G218gat), .B1(new_n930_), .B2(new_n646_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1355gat));
endmodule


