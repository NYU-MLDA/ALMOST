//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT70), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n210_));
  AND3_X1   g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n206_), .B2(new_n209_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214_));
  INV_X1    g013(.A(G1gat), .ZN(new_n215_));
  INV_X1    g014(.A(G8gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n217_), .B2(KEYINPUT74), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(KEYINPUT74), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G1gat), .B(G8gat), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n206_), .A2(new_n209_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n224_), .B(new_n225_), .C1(new_n223_), .C2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n225_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n223_), .A2(new_n226_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n223_), .A2(new_n226_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G169gat), .B(G197gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(G43gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT78), .B(G15gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT23), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT76), .B(G183gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(G190gat), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G169gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n248_), .B(KEYINPUT23), .ZN(new_n255_));
  OR3_X1    g054(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT26), .B(G190gat), .Z(new_n258_));
  NOR2_X1   g057(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(new_n250_), .B2(KEYINPUT25), .ZN(new_n260_));
  OAI22_X1  g059(.A1(new_n257_), .A2(KEYINPUT77), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G169gat), .ZN(new_n264_));
  INV_X1    g063(.A(G176gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n255_), .A2(new_n256_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT77), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n254_), .B1(new_n261_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT30), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT79), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n247_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n273_), .B2(new_n247_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G127gat), .B(G134gat), .Z(new_n277_));
  XOR2_X1   g076(.A(G113gat), .B(G120gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n279_), .B(KEYINPUT31), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n276_), .A2(new_n281_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT85), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G155gat), .B(G162gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT2), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n289_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n289_), .A2(KEYINPUT1), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n291_), .A2(new_n292_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n294_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT29), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT82), .B(G204gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(G197gat), .ZN(new_n311_));
  INV_X1    g110(.A(G197gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(G204gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT21), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G197gat), .A2(G204gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n314_), .B(new_n315_), .C1(new_n319_), .C2(KEYINPUT21), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n315_), .B(KEYINPUT83), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(KEYINPUT84), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n323_), .B(new_n317_), .C1(new_n310_), .C2(new_n312_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n321_), .A2(new_n322_), .A3(KEYINPUT21), .A4(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(G228gat), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n309_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n309_), .B2(new_n326_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n288_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT86), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n308_), .A2(KEYINPUT29), .ZN(new_n335_));
  XOR2_X1   g134(.A(G22gat), .B(G50gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT28), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n331_), .A2(new_n332_), .A3(new_n288_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n333_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n334_), .A2(new_n338_), .B1(new_n340_), .B2(new_n333_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n279_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n308_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n302_), .A2(new_n307_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n279_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT91), .Z(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G85gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT0), .B(G57gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT93), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(new_n360_), .A3(new_n357_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n347_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n348_), .A2(KEYINPUT4), .A3(new_n279_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n350_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n351_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n366_), .A2(KEYINPUT33), .A3(new_n367_), .A4(new_n356_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n356_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT92), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n374_), .A3(new_n371_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n369_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n326_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT25), .B(G183gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT88), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n266_), .B(new_n257_), .C1(new_n384_), .C2(new_n258_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n249_), .B1(G183gat), .B2(G190gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n253_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n382_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT19), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT20), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n270_), .B2(new_n326_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT89), .B1(new_n326_), .B2(new_n388_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n391_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n393_), .B(KEYINPUT87), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n270_), .A2(new_n326_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n326_), .B2(new_n388_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n381_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n403_), .B1(new_n326_), .B2(new_n270_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n399_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n397_), .A3(new_n380_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n405_), .A2(new_n408_), .A3(KEYINPUT90), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT90), .B1(new_n405_), .B2(new_n408_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n376_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n398_), .A2(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT94), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT95), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(KEYINPUT95), .A3(new_n414_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n366_), .A2(new_n367_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n357_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n370_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n406_), .A2(new_n399_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n382_), .A2(new_n389_), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n270_), .B2(new_n326_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n393_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT32), .B(new_n380_), .C1(new_n422_), .C2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n417_), .A2(new_n418_), .A3(new_n421_), .A4(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n345_), .B1(new_n411_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n405_), .A2(new_n408_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n381_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(KEYINPUT27), .A3(new_n408_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n435_), .A2(new_n344_), .A3(new_n421_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n285_), .B1(new_n429_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n344_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT97), .ZN(new_n439_));
  INV_X1    g238(.A(new_n421_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n344_), .A2(new_n441_), .A3(new_n432_), .A4(new_n434_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n439_), .A2(new_n284_), .A3(new_n440_), .A4(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n240_), .B1(new_n437_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G190gat), .B(G218gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G134gat), .B(G162gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(KEYINPUT36), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT68), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT65), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT65), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n454_));
  AND2_X1   g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G85gat), .ZN(new_n463_));
  INV_X1    g262(.A(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT9), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT64), .B(G85gat), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n464_), .A2(KEYINPUT9), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n462_), .B(new_n467_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n450_), .B1(new_n458_), .B2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n462_), .A2(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n451_), .A2(KEYINPUT65), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n468_), .A2(new_n469_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n472_), .A2(new_n478_), .A3(new_n479_), .A4(KEYINPUT68), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  INV_X1    g280(.A(G99gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n460_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n465_), .A2(new_n466_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n486_), .A2(KEYINPUT8), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT8), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n483_), .A2(new_n484_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n487_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n471_), .B(new_n480_), .C1(new_n488_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n213_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT34), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT72), .B1(new_n497_), .B2(KEYINPUT35), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n458_), .A2(new_n470_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT8), .B1(new_n486_), .B2(new_n487_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n491_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n226_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n498_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n495_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n495_), .A2(new_n506_), .A3(new_n504_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n449_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n447_), .A2(KEYINPUT36), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n511_), .A3(new_n509_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT73), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n508_), .A2(KEYINPUT73), .A3(new_n511_), .A4(new_n509_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n510_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G176gat), .B(G204gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  NAND2_X1  g321(.A1(G230gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G78gat), .Z(new_n526_));
  OR2_X1    g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n472_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n530_), .B(new_n531_), .C1(new_n488_), .C2(new_n493_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT66), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n502_), .A2(KEYINPUT66), .A3(new_n530_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT67), .A3(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n502_), .A2(new_n530_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT67), .B1(new_n534_), .B2(new_n535_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n523_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n502_), .B2(new_n530_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n523_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n502_), .B2(new_n530_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n527_), .B(KEYINPUT12), .C1(new_n529_), .C2(new_n528_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n488_), .A2(new_n493_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n471_), .A2(new_n480_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n543_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n543_), .A2(new_n545_), .A3(new_n550_), .A4(KEYINPUT69), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n522_), .B1(new_n541_), .B2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n553_), .A2(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n536_), .A2(new_n537_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n544_), .B1(new_n558_), .B2(new_n539_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n522_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n561_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT75), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n223_), .B(new_n567_), .Z(new_n568_));
  AND2_X1   g367(.A1(new_n568_), .A2(new_n530_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n530_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT17), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  OAI211_X1 g377(.A(KEYINPUT17), .B(new_n578_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n566_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT75), .B1(new_n571_), .B2(new_n576_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n518_), .A2(new_n562_), .A3(new_n565_), .A4(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n444_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT98), .Z(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n215_), .A3(new_n421_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n516_), .B1(new_n437_), .B2(new_n443_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n565_), .A2(new_n562_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n239_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n582_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n215_), .B1(new_n596_), .B2(new_n421_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n589_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n588_), .B2(new_n587_), .ZN(G1324gat));
  NAND3_X1  g398(.A1(new_n586_), .A2(new_n216_), .A3(new_n435_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n435_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G8gat), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT39), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(KEYINPUT39), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(G1325gat));
  OR3_X1    g406(.A1(new_n585_), .A2(G15gat), .A3(new_n285_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n596_), .A2(new_n284_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT41), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(G15gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n609_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n612_), .B1(new_n611_), .B2(G15gat), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1326gat));
  OR3_X1    g419(.A1(new_n585_), .A2(G22gat), .A3(new_n344_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n596_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G22gat), .B1(new_n622_), .B2(new_n344_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(KEYINPUT42), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(KEYINPUT42), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1327gat));
  NAND2_X1  g427(.A1(new_n514_), .A2(new_n515_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n510_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n582_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n591_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n444_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n421_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n593_), .A2(new_n582_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n437_), .A2(new_n443_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n516_), .B(KEYINPUT37), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  AOI211_X1 g441(.A(KEYINPUT43), .B(new_n518_), .C1(new_n437_), .C2(new_n443_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT44), .B(new_n638_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n421_), .A2(G29gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n637_), .B1(new_n648_), .B2(new_n649_), .ZN(G1328gat));
  XNOR2_X1  g449(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(new_n435_), .A3(new_n647_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G36gat), .ZN(new_n653_));
  INV_X1    g452(.A(G36gat), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n444_), .A2(new_n654_), .A3(new_n435_), .A4(new_n634_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n653_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n651_), .B1(new_n659_), .B2(KEYINPUT103), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n652_), .B2(G36gat), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662_));
  INV_X1    g461(.A(new_n651_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n660_), .A2(new_n664_), .ZN(G1329gat));
  NAND4_X1  g464(.A1(new_n646_), .A2(G43gat), .A3(new_n284_), .A4(new_n647_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n242_), .B1(new_n635_), .B2(new_n285_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g468(.A1(new_n646_), .A2(new_n345_), .A3(new_n647_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G50gat), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n635_), .A2(G50gat), .A3(new_n344_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT105), .ZN(G1331gat));
  AOI21_X1  g473(.A(new_n239_), .B1(new_n437_), .B2(new_n443_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n641_), .A2(new_n594_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(new_n591_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(G57gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n421_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n592_), .A2(new_n239_), .A3(new_n594_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n590_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n440_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1332gat));
  INV_X1    g482(.A(G64gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n681_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n435_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT48), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n677_), .A2(new_n684_), .A3(new_n435_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1333gat));
  INV_X1    g488(.A(G71gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n677_), .A2(new_n690_), .A3(new_n284_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G71gat), .B1(new_n681_), .B2(new_n285_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT49), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT49), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT106), .Z(G1334gat));
  OAI21_X1  g495(.A(G78gat), .B1(new_n681_), .B2(new_n344_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT50), .ZN(new_n698_));
  INV_X1    g497(.A(G78gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n677_), .A2(new_n699_), .A3(new_n345_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1335gat));
  OR2_X1    g500(.A1(new_n642_), .A2(new_n643_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n592_), .A2(new_n239_), .A3(new_n582_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n440_), .A2(new_n468_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n633_), .A2(new_n592_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n675_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n463_), .B1(new_n708_), .B2(new_n440_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT107), .ZN(G1336gat));
  INV_X1    g510(.A(new_n708_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G92gat), .B1(new_n712_), .B2(new_n435_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT108), .Z(new_n714_));
  AOI21_X1  g513(.A(new_n464_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n704_), .B2(new_n715_), .ZN(G1337gat));
  NAND4_X1  g515(.A1(new_n712_), .A2(new_n284_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n284_), .B(new_n703_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT109), .B1(new_n718_), .B2(G99gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n712_), .A2(new_n460_), .A3(new_n345_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n345_), .B(new_n703_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(new_n725_), .A3(G106gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n724_), .B2(G106gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g528(.A(KEYINPUT59), .ZN(new_n730_));
  XOR2_X1   g529(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n583_), .B2(new_n239_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n676_), .A2(new_n240_), .A3(new_n592_), .A4(new_n731_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(KEYINPUT112), .A2(KEYINPUT56), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n551_), .A2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n543_), .A2(new_n550_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n532_), .A2(new_n533_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT66), .B1(new_n502_), .B2(new_n530_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(new_n743_), .A3(KEYINPUT111), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n543_), .A2(new_n534_), .A3(new_n550_), .A4(new_n535_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n739_), .B1(new_n748_), .B2(new_n544_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n553_), .A2(new_n738_), .A3(new_n554_), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n560_), .B(new_n737_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT111), .B1(new_n740_), .B2(new_n743_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n745_), .A2(new_n746_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n544_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n739_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n750_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n736_), .B1(new_n756_), .B2(new_n522_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n239_), .A2(new_n561_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n751_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n230_), .A2(new_n225_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n224_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n225_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n236_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT113), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n224_), .A2(new_n760_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n236_), .A4(new_n762_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n238_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n560_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n563_), .A2(new_n774_), .A3(new_n769_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n631_), .B1(new_n759_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT57), .B(new_n631_), .C1(new_n759_), .C2(new_n776_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n770_), .A2(new_n768_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n560_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n756_), .A2(new_n784_), .A3(new_n522_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n781_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n523_), .B1(new_n744_), .B2(new_n747_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n553_), .A2(new_n738_), .A3(new_n554_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n739_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n560_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT58), .A3(new_n786_), .A4(new_n782_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n788_), .A2(new_n641_), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n779_), .A2(new_n780_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n735_), .B1(new_n795_), .B2(new_n594_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n730_), .B1(new_n796_), .B2(KEYINPUT115), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n439_), .A2(new_n284_), .A3(new_n442_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n793_), .A2(new_n641_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n778_), .A2(new_n777_), .B1(new_n799_), .B2(new_n788_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n582_), .B1(new_n800_), .B2(new_n780_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n421_), .B(new_n798_), .C1(new_n801_), .C2(new_n735_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n797_), .B(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n240_), .ZN(new_n804_));
  OR3_X1    g603(.A1(new_n802_), .A2(G113gat), .A3(new_n240_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1340gat));
  INV_X1    g605(.A(new_n803_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n802_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT60), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT116), .B(G120gat), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n592_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n592_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n808_), .A2(new_n809_), .A3(new_n812_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n807_), .A2(new_n813_), .B1(new_n814_), .B2(new_n810_), .ZN(G1341gat));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n802_), .B2(new_n594_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n594_), .A2(new_n819_), .A3(new_n817_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n819_), .B2(new_n817_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n816_), .B(new_n818_), .C1(new_n803_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n801_), .B2(new_n735_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n802_), .A2(new_n730_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n774_), .B1(new_n563_), .B2(new_n769_), .ZN(new_n826_));
  AOI211_X1 g625(.A(KEYINPUT114), .B(new_n768_), .C1(new_n556_), .C2(new_n561_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n756_), .A2(new_n522_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n737_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n783_), .A2(new_n736_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n758_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n516_), .B1(new_n828_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n794_), .B1(new_n834_), .B2(KEYINPUT57), .ZN(new_n835_));
  INV_X1    g634(.A(new_n780_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n594_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n735_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n440_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT115), .B1(new_n837_), .B2(new_n838_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n798_), .B(new_n839_), .C1(new_n840_), .C2(KEYINPUT59), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n821_), .B1(new_n825_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n818_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n822_), .A2(new_n844_), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n802_), .B2(new_n631_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n641_), .A2(G134gat), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT119), .B(new_n847_), .C1(new_n803_), .C2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n825_), .B2(new_n841_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n847_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n285_), .A2(new_n345_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n435_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n839_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n239_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n591_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g660(.A1(new_n839_), .A2(new_n582_), .A3(new_n856_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n862_), .A2(KEYINPUT120), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(KEYINPUT120), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1346gat));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n857_), .A2(new_n869_), .A3(new_n516_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n857_), .A2(new_n641_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1347gat));
  NAND2_X1  g671(.A1(new_n837_), .A2(new_n838_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT22), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n435_), .A2(new_n440_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n285_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n239_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n873_), .A2(new_n874_), .A3(new_n344_), .A4(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(KEYINPUT62), .A3(new_n264_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n796_), .A2(new_n345_), .A3(new_n877_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n874_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n873_), .A2(new_n881_), .A3(new_n344_), .A4(new_n878_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G169gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n880_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT121), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n888_), .B(new_n880_), .C1(new_n883_), .C2(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1348gat));
  NOR2_X1   g689(.A1(new_n796_), .A2(new_n345_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n876_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n592_), .B1(KEYINPUT122), .B2(new_n265_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n265_), .A2(KEYINPUT122), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1349gat));
  NOR2_X1   g696(.A1(new_n892_), .A2(new_n594_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n250_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n384_), .B2(new_n898_), .ZN(G1350gat));
  OR3_X1    g699(.A1(new_n892_), .A2(new_n258_), .A3(new_n631_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n891_), .A2(new_n641_), .A3(new_n876_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n902_), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT123), .B1(new_n902_), .B2(G190gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n901_), .B1(new_n903_), .B2(new_n904_), .ZN(G1351gat));
  NOR3_X1   g704(.A1(new_n796_), .A2(new_n855_), .A3(new_n875_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G197gat), .B1(new_n906_), .B2(new_n239_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n907_), .A2(KEYINPUT125), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(KEYINPUT125), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n906_), .A2(G197gat), .A3(new_n239_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n910_), .A2(KEYINPUT124), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(KEYINPUT124), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n908_), .A2(new_n909_), .B1(new_n911_), .B2(new_n912_), .ZN(G1352gat));
  INV_X1    g712(.A(G204gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n906_), .B2(new_n591_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n906_), .A2(new_n310_), .A3(new_n591_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n916_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(G1353gat));
  NOR2_X1   g719(.A1(new_n855_), .A2(new_n875_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n873_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n594_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AND2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n923_), .B2(new_n924_), .ZN(G1354gat));
  AND3_X1   g726(.A1(new_n906_), .A2(G218gat), .A3(new_n641_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n922_), .A2(new_n631_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n929_), .A2(KEYINPUT127), .ZN(new_n930_));
  AOI21_X1  g729(.A(G218gat), .B1(new_n929_), .B2(KEYINPUT127), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n930_), .B2(new_n931_), .ZN(G1355gat));
endmodule


