//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n207_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NOR4_X1   g015(.A1(KEYINPUT88), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(G141gat), .B2(G148gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n206_), .A2(KEYINPUT2), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n223_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT89), .B1(new_n222_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT88), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n219_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n206_), .A2(KEYINPUT2), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n224_), .A2(G141gat), .A3(G148gat), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n234_), .A2(new_n235_), .B1(new_n205_), .B2(KEYINPUT3), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n228_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n214_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n216_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT29), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n202_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(new_n228_), .B2(new_n237_), .ZN(new_n244_));
  NOR4_X1   g043(.A1(new_n244_), .A2(KEYINPUT28), .A3(new_n216_), .A4(KEYINPUT29), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT90), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G22gat), .B(G50gat), .Z(new_n247_));
  AND3_X1   g046(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n233_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n239_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n216_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n241_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT28), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n240_), .A2(new_n202_), .A3(new_n241_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT90), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n246_), .A2(new_n247_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n247_), .B1(new_n246_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT29), .B1(new_n244_), .B2(new_n216_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT93), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262_));
  INV_X1    g061(.A(G197gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT91), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G197gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n262_), .B1(new_n267_), .B2(G204gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n261_), .B1(new_n268_), .B2(KEYINPUT21), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT92), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n263_), .B2(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT91), .B(G197gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(G204gat), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n267_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n275_), .A3(KEYINPUT21), .ZN(new_n276_));
  INV_X1    g075(.A(new_n262_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT21), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(KEYINPUT93), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT94), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT94), .ZN(new_n283_));
  INV_X1    g082(.A(G211gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n284_), .A2(G218gat), .ZN(new_n285_));
  INV_X1    g084(.A(G218gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(G211gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n283_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n282_), .A2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n269_), .A2(new_n276_), .A3(new_n280_), .A4(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT95), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n282_), .A2(new_n288_), .A3(KEYINPUT95), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT21), .A4(new_n268_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n260_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n260_), .A2(new_n297_), .A3(new_n295_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G78gat), .B(G106gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n302_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n259_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n260_), .A2(new_n297_), .A3(new_n295_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n297_), .B1(new_n260_), .B2(new_n295_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT96), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT96), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n299_), .A2(new_n310_), .A3(new_n300_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n311_), .A3(new_n302_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT97), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT97), .A4(new_n302_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n314_), .A2(new_n259_), .A3(new_n304_), .A4(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT98), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n257_), .A2(new_n303_), .A3(new_n258_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(KEYINPUT98), .A3(new_n315_), .A4(new_n314_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n306_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G71gat), .B(G99gat), .ZN(new_n322_));
  INV_X1    g121(.A(G43gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT30), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(G15gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n325_), .A2(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT83), .ZN(new_n334_));
  INV_X1    g133(.A(G183gat), .ZN(new_n335_));
  INV_X1    g134(.A(G190gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT23), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n334_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(KEYINPUT26), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n339_), .A2(KEYINPUT82), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n336_), .A2(KEYINPUT26), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(KEYINPUT82), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(KEYINPUT24), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n349_), .B2(KEYINPUT24), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n338_), .A2(new_n344_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n337_), .A2(new_n333_), .A3(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n332_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n353_), .B(new_n354_), .C1(G183gat), .C2(G190gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G169gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n351_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT86), .B1(new_n331_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT31), .ZN(new_n364_));
  XOR2_X1   g163(.A(G127gat), .B(G134gat), .Z(new_n365_));
  INV_X1    g164(.A(KEYINPUT85), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT85), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G113gat), .B(G120gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n364_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT104), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT103), .B(KEYINPUT18), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n380_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT20), .B1(new_n295_), .B2(new_n359_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT100), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT100), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT24), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n389_), .A3(new_n345_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n353_), .A2(new_n354_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT101), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT101), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n353_), .A2(new_n393_), .A3(new_n354_), .A4(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n342_), .B(KEYINPUT99), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n341_), .A2(new_n339_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n387_), .A2(new_n389_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n396_), .A2(new_n397_), .B1(new_n398_), .B2(new_n349_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n338_), .B1(G183gat), .B2(G190gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n348_), .B(KEYINPUT102), .ZN(new_n402_));
  INV_X1    g201(.A(G176gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT22), .B(G169gat), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n400_), .A2(new_n406_), .B1(new_n294_), .B2(new_n290_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT19), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n385_), .A2(new_n408_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n295_), .B2(new_n359_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n400_), .A2(new_n406_), .A3(new_n294_), .A4(new_n290_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n410_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n383_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n410_), .B1(new_n384_), .B2(new_n407_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n419_), .A2(new_n383_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  OR3_X1    g221(.A1(new_n418_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n383_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n374_), .B1(new_n244_), .B2(new_n216_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n367_), .A2(new_n369_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n370_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n371_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n250_), .A2(new_n432_), .A3(new_n251_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n433_), .A3(KEYINPUT4), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n374_), .B(new_n435_), .C1(new_n244_), .C2(new_n216_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n437_), .B(KEYINPUT105), .Z(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n428_), .A2(new_n433_), .A3(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT106), .B(G85gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT0), .B(G57gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT108), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n439_), .A2(new_n440_), .A3(new_n446_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n441_), .A2(KEYINPUT108), .A3(new_n447_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n321_), .A2(new_n375_), .A3(new_n427_), .A4(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n364_), .B(new_n432_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n453_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n426_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n321_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n318_), .A2(new_n320_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n306_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n450_), .A2(KEYINPUT107), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT33), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n421_), .A2(new_n424_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n450_), .A2(KEYINPUT107), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n434_), .A2(new_n437_), .A3(new_n436_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n428_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n447_), .A3(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .A4(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n381_), .A2(KEYINPUT32), .A3(new_n382_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n419_), .A2(new_n420_), .A3(new_n470_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n459_), .A2(new_n460_), .A3(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n454_), .B1(new_n458_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G169gat), .B(G197gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT80), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G113gat), .B(G141gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485_));
  INV_X1    g284(.A(G1gat), .ZN(new_n486_));
  INV_X1    g285(.A(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G8gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G29gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n491_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n494_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n491_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n491_), .A2(new_n495_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n497_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n484_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506_));
  INV_X1    g305(.A(new_n504_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n499_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n483_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n483_), .B(KEYINPUT81), .C1(new_n507_), .C2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n477_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT109), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G85gat), .B(G92gat), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT9), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT6), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(G99gat), .A3(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G85gat), .ZN(new_n526_));
  INV_X1    g325(.A(G92gat), .ZN(new_n527_));
  OR3_X1    g326(.A1(new_n526_), .A2(new_n527_), .A3(KEYINPUT9), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n518_), .A2(new_n520_), .A3(new_n525_), .A4(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT8), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n522_), .A2(new_n524_), .A3(KEYINPUT65), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n537_));
  OAI22_X1  g336(.A1(new_n536_), .A2(new_n537_), .B1(G99gat), .B2(G106gat), .ZN(new_n538_));
  INV_X1    g337(.A(G99gat), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n517_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n532_), .A2(new_n533_), .A3(new_n538_), .A4(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n530_), .B1(new_n541_), .B2(new_n519_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n519_), .A2(new_n530_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n538_), .A2(new_n540_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n525_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n529_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n549_));
  XOR2_X1   g348(.A(G71gat), .B(G78gat), .Z(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT66), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT12), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT66), .B1(new_n546_), .B2(new_n554_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n546_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n553_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n558_), .A2(new_n559_), .A3(new_n562_), .A4(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n555_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n559_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G120gat), .B(G148gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(G176gat), .B(G204gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n565_), .A2(new_n568_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n565_), .A2(new_n568_), .A3(KEYINPUT70), .A4(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n565_), .A2(new_n568_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT67), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n565_), .A2(new_n568_), .A3(KEYINPUT67), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n573_), .B(KEYINPUT69), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n578_), .A2(new_n584_), .A3(KEYINPUT13), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT13), .B1(new_n578_), .B2(new_n584_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n491_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n553_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT76), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(KEYINPUT76), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n593_), .A2(new_n594_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n591_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n563_), .A2(new_n494_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n546_), .A2(new_n501_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n610_), .A2(new_n611_), .A3(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n615_), .A2(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n621_));
  INV_X1    g420(.A(new_n619_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n610_), .A2(new_n611_), .A3(new_n622_), .A4(new_n617_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n621_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n609_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n624_), .B2(KEYINPUT73), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n629_), .B(new_n609_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n605_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n588_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n515_), .A2(new_n486_), .A3(new_n456_), .A4(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n635_), .A2(KEYINPUT110), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n459_), .A2(new_n460_), .A3(new_n475_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(new_n455_), .C1(new_n321_), .C2(new_n457_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n627_), .B1(new_n639_), .B2(new_n454_), .ZN(new_n640_));
  NOR4_X1   g439(.A1(new_n586_), .A2(new_n587_), .A3(new_n512_), .A4(new_n605_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n486_), .B1(new_n642_), .B2(new_n456_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n635_), .B1(new_n636_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT110), .B1(new_n635_), .B2(new_n636_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n644_), .A3(new_n645_), .ZN(G1324gat));
  XNOR2_X1  g445(.A(KEYINPUT112), .B(KEYINPUT39), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n640_), .A2(KEYINPUT111), .A3(new_n426_), .A4(new_n641_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n627_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n477_), .A2(new_n426_), .A3(new_n650_), .A4(new_n641_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT111), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n647_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n654_));
  AND4_X1   g453(.A1(G8gat), .A2(new_n653_), .A3(new_n648_), .A4(new_n647_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n515_), .A2(new_n634_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n426_), .A2(new_n487_), .ZN(new_n657_));
  OAI22_X1  g456(.A1(new_n654_), .A2(new_n655_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI221_X1 g459(.A(KEYINPUT40), .B1(new_n656_), .B2(new_n657_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  INV_X1    g461(.A(KEYINPUT113), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n375_), .A2(new_n327_), .ZN(new_n664_));
  OR3_X1    g463(.A1(new_n656_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n327_), .B1(new_n642_), .B2(new_n375_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT41), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n656_), .B2(new_n664_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n667_), .A3(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n321_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n642_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT42), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n670_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n656_), .B2(new_n674_), .ZN(G1327gat));
  INV_X1    g474(.A(new_n605_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n650_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n588_), .A2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n515_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n456_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n588_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(new_n512_), .A3(new_n676_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n631_), .A2(new_n632_), .ZN(new_n683_));
  AND2_X1   g482(.A1(KEYINPUT114), .A2(KEYINPUT43), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n683_), .B(new_n684_), .C1(new_n639_), .C2(new_n454_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(KEYINPUT114), .A2(KEYINPUT43), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n683_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n477_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n682_), .B1(new_n685_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n682_), .C1(new_n685_), .C2(new_n689_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n456_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n680_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n692_), .A2(new_n426_), .A3(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n427_), .A2(G36gat), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n515_), .A2(new_n699_), .A3(new_n678_), .A4(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n514_), .A2(KEYINPUT109), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n477_), .B2(new_n513_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n678_), .B(new_n700_), .C1(new_n702_), .C2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT45), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n698_), .A2(KEYINPUT46), .A3(new_n707_), .ZN(new_n708_));
  AOI22_X1  g507(.A1(new_n697_), .A2(G36gat), .B1(new_n701_), .B2(new_n706_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT115), .B(KEYINPUT46), .Z(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(G1329gat));
  NAND3_X1  g510(.A1(new_n515_), .A2(new_n375_), .A3(new_n678_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n323_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n692_), .A2(G43gat), .A3(new_n375_), .A4(new_n693_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT47), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1330gat));
  INV_X1    g518(.A(G50gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n679_), .A2(new_n720_), .A3(new_n671_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT116), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n694_), .B2(new_n671_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n692_), .A2(new_n722_), .A3(new_n671_), .A4(new_n693_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G50gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n723_), .B2(new_n725_), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n588_), .A2(new_n513_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n640_), .A2(new_n676_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n453_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n477_), .A2(new_n727_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n633_), .ZN(new_n732_));
  INV_X1    g531(.A(G57gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n456_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1332gat));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n728_), .B2(new_n426_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT48), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n732_), .A2(new_n736_), .A3(new_n426_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n728_), .B2(new_n375_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT49), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n732_), .A2(new_n741_), .A3(new_n375_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1334gat));
  INV_X1    g544(.A(G78gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n732_), .A2(new_n746_), .A3(new_n671_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n728_), .A2(new_n671_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G78gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT50), .B(new_n746_), .C1(new_n728_), .C2(new_n671_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT117), .B(new_n747_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1335gat));
  AND2_X1   g555(.A1(new_n731_), .A2(new_n677_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n526_), .A3(new_n456_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n685_), .A2(new_n689_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n727_), .A2(new_n605_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n759_), .A2(new_n453_), .A3(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n761_), .B2(new_n526_), .ZN(G1336gat));
  NAND3_X1  g561(.A1(new_n757_), .A2(new_n527_), .A3(new_n426_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n759_), .A2(new_n427_), .A3(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n527_), .ZN(G1337gat));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n375_), .A2(new_n516_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n757_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n760_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n375_), .B(new_n769_), .C1(new_n685_), .C2(new_n689_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(KEYINPUT118), .A3(G99gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT118), .B1(new_n770_), .B2(G99gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n768_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n757_), .A2(new_n517_), .A3(new_n671_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n671_), .B(new_n769_), .C1(new_n685_), .C2(new_n689_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n778_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NOR4_X1   g586(.A1(new_n671_), .A2(new_n426_), .A3(new_n455_), .A4(new_n453_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n578_), .A2(new_n584_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n502_), .A2(new_n503_), .A3(new_n498_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n496_), .A2(new_n497_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n483_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n505_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n583_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n562_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n564_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n567_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT55), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n565_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NOR4_X1   g600(.A1(new_n796_), .A2(new_n797_), .A3(new_n801_), .A4(new_n567_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n795_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n512_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n794_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n650_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n796_), .A2(new_n797_), .A3(new_n567_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(KEYINPUT55), .B2(new_n798_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n583_), .B1(new_n814_), .B2(new_n802_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT56), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n804_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n505_), .A2(new_n793_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n683_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n816_), .A2(new_n818_), .A3(KEYINPUT58), .A4(new_n820_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n811_), .A2(new_n812_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n810_), .A2(KEYINPUT57), .A3(new_n650_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n676_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n587_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(new_n633_), .A3(new_n512_), .A4(new_n585_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n831_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n588_), .A2(new_n512_), .A3(new_n633_), .A4(new_n833_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n832_), .A2(new_n834_), .B1(KEYINPUT120), .B2(KEYINPUT54), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n788_), .B(new_n789_), .C1(new_n827_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT123), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n811_), .A2(new_n812_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n823_), .A2(new_n824_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n826_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n605_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n835_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n788_), .A4(new_n789_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n835_), .B1(new_n840_), .B2(new_n605_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n788_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT59), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n837_), .A2(new_n845_), .A3(new_n513_), .A4(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G113gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n843_), .A2(new_n788_), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n851_), .A2(G113gat), .A3(new_n512_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1340gat));
  NAND4_X1  g652(.A1(new_n837_), .A2(new_n845_), .A3(new_n681_), .A4(new_n848_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT124), .B(G120gat), .Z(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n855_), .A2(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n588_), .B2(KEYINPUT60), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n843_), .A2(new_n788_), .A3(new_n858_), .A4(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n862_), .ZN(G1341gat));
  NAND4_X1  g662(.A1(new_n837_), .A2(new_n845_), .A3(new_n676_), .A4(new_n848_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G127gat), .ZN(new_n865_));
  OR3_X1    g664(.A1(new_n851_), .A2(G127gat), .A3(new_n605_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1342gat));
  NAND4_X1  g666(.A1(new_n837_), .A2(new_n845_), .A3(new_n688_), .A4(new_n848_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G134gat), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n851_), .A2(G134gat), .A3(new_n650_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1343gat));
  NOR3_X1   g670(.A1(new_n846_), .A2(new_n321_), .A3(new_n375_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n426_), .A2(new_n453_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n203_), .A3(new_n513_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n873_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G141gat), .B1(new_n876_), .B2(new_n512_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n204_), .A3(new_n681_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G148gat), .B1(new_n876_), .B2(new_n588_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1345gat));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n874_), .A2(new_n676_), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n876_), .B2(new_n605_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n876_), .B2(new_n683_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n650_), .A2(G162gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n876_), .B2(new_n888_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n846_), .A2(new_n671_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n455_), .A2(new_n427_), .A3(new_n456_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n404_), .A3(new_n513_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n843_), .A2(new_n321_), .A3(new_n513_), .A4(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G169gat), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(new_n898_), .A3(new_n899_), .ZN(G1348gat));
  OAI21_X1  g699(.A(new_n403_), .B1(new_n892_), .B2(new_n588_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n846_), .B2(new_n671_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n681_), .A2(G176gat), .A3(new_n891_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n901_), .A2(new_n906_), .ZN(G1349gat));
  OR2_X1    g706(.A1(new_n605_), .A2(new_n396_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n892_), .A2(new_n908_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n902_), .A2(new_n676_), .A3(new_n891_), .A4(new_n904_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n335_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n892_), .B2(new_n683_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n627_), .A2(new_n397_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n892_), .B2(new_n913_), .ZN(G1351gat));
  NOR2_X1   g713(.A1(new_n427_), .A2(new_n456_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n872_), .A2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT127), .B(G197gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n513_), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n917_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n872_), .A2(new_n915_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n512_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n921_), .ZN(G1352gat));
  NAND3_X1  g721(.A1(new_n916_), .A2(new_n274_), .A3(new_n681_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G204gat), .B1(new_n920_), .B2(new_n588_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1353gat));
  NOR2_X1   g724(.A1(new_n321_), .A2(new_n375_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n843_), .A2(new_n676_), .A3(new_n926_), .A4(new_n915_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  AND2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n927_), .B2(new_n928_), .ZN(G1354gat));
  NAND3_X1  g730(.A1(new_n916_), .A2(new_n286_), .A3(new_n627_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G218gat), .B1(new_n920_), .B2(new_n683_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1355gat));
endmodule


