//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT31), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207_));
  INV_X1    g006(.A(G15gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT79), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G71gat), .B(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G43gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n210_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT22), .ZN(new_n215_));
  OR2_X1    g014(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT78), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT78), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(new_n215_), .B2(G169gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n219_), .B(new_n220_), .C1(new_n218_), .C2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT23), .ZN(new_n227_));
  OR2_X1    g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n225_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G169gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n220_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT25), .B(G183gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT26), .B(G190gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n223_), .A2(new_n229_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n238_), .A2(KEYINPUT30), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(KEYINPUT30), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n214_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT80), .B(new_n214_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n239_), .A2(new_n240_), .A3(new_n214_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n206_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  AOI211_X1 g047(.A(KEYINPUT31), .B(new_n246_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n205_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n244_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n238_), .B(KEYINPUT30), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT80), .B1(new_n252_), .B2(new_n214_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n247_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT31), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n245_), .A2(new_n206_), .A3(new_n247_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n204_), .A3(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT83), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n259_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n260_), .B1(KEYINPUT83), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT2), .ZN(new_n264_));
  OR2_X1    g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n259_), .A3(KEYINPUT3), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n269_), .B2(KEYINPUT1), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(KEYINPUT82), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n272_), .A2(KEYINPUT82), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n263_), .B(new_n265_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n204_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n204_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(KEYINPUT4), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n277_), .A2(new_n205_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(new_n280_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G1gat), .B(G29gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n286_), .A2(new_n289_), .A3(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n258_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT100), .ZN(new_n302_));
  INV_X1    g101(.A(G233gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n303_), .A2(KEYINPUT84), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(KEYINPUT84), .ZN(new_n305_));
  OAI21_X1  g104(.A(G228gat), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n309_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n309_), .B2(new_n315_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n306_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT87), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n309_), .A2(new_n315_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n312_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n309_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n322_), .A2(new_n326_), .A3(new_n327_), .A4(new_n306_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n326_), .B1(new_n278_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n306_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n321_), .A2(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(KEYINPUT89), .A3(new_n334_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT89), .B1(new_n332_), .B2(new_n334_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n336_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n277_), .A2(KEYINPUT29), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G22gat), .B(G50gat), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n343_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n340_), .A2(KEYINPUT90), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT90), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n321_), .A2(new_n328_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n330_), .A2(new_n331_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n334_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n335_), .B1(new_n354_), .B2(new_n337_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n349_), .B1(new_n355_), .B2(new_n346_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n351_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT91), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n333_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT91), .B1(new_n332_), .B2(new_n334_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n346_), .A2(new_n359_), .A3(new_n352_), .A4(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n348_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT27), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n316_), .A2(new_n317_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT95), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n220_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n225_), .A2(KEYINPUT94), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n225_), .A2(KEYINPUT94), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n228_), .A2(new_n227_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n227_), .A2(new_n232_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(new_n234_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT93), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n236_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n236_), .A2(new_n377_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n235_), .A3(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n371_), .A2(new_n374_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n367_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n223_), .A2(new_n229_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n233_), .A2(new_n237_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT20), .B1(new_n326_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT92), .B(KEYINPUT20), .C1(new_n326_), .C2(new_n385_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n366_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n367_), .B2(new_n381_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n367_), .A2(KEYINPUT96), .A3(new_n238_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT96), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n326_), .B2(new_n385_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n366_), .B(new_n392_), .C1(new_n393_), .C2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n390_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT18), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  AOI21_X1  g201(.A(new_n363_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT99), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n371_), .A2(new_n374_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n376_), .A2(new_n380_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n324_), .A2(new_n405_), .A3(new_n325_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT20), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT96), .B1(new_n367_), .B2(new_n238_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n326_), .A2(new_n385_), .A3(new_n394_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n404_), .B1(new_n411_), .B2(new_n366_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n388_), .A2(new_n366_), .A3(new_n389_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n392_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(KEYINPUT99), .A3(new_n365_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n402_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n403_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n417_), .B1(new_n390_), .B2(new_n397_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n386_), .A2(new_n387_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n382_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n389_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n365_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n402_), .A3(new_n396_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n363_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n419_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n302_), .B1(new_n362_), .B2(new_n428_), .ZN(new_n429_));
  AND4_X1   g228(.A1(new_n346_), .A2(new_n359_), .A3(new_n360_), .A4(new_n352_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n354_), .A2(new_n337_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n346_), .B1(new_n431_), .B2(new_n336_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n432_), .B2(KEYINPUT90), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n418_), .A2(new_n403_), .B1(new_n426_), .B2(new_n363_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(KEYINPUT100), .A4(new_n356_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n301_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n250_), .A2(new_n257_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n362_), .A2(new_n300_), .A3(new_n434_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n402_), .A2(KEYINPUT32), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n416_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n424_), .A2(new_n396_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n299_), .B1(new_n445_), .B2(new_n443_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n286_), .A2(new_n289_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT33), .A4(new_n295_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n282_), .B(new_n283_), .C1(KEYINPUT4), .C2(new_n281_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n283_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n295_), .B1(new_n288_), .B2(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n298_), .A2(new_n450_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT98), .B1(new_n298_), .B2(new_n450_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n449_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  OAI22_X1  g255(.A1(new_n444_), .A2(new_n446_), .B1(new_n456_), .B2(new_n426_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n433_), .A3(new_n356_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n440_), .B1(new_n441_), .B2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n436_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G8gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G43gat), .B(G50gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n467_), .B(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n473_), .A2(G229gat), .A3(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n475_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n467_), .A2(new_n472_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n472_), .B(KEYINPUT15), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n480_), .B2(new_n467_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n476_), .A2(new_n477_), .A3(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G169gat), .B(G197gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT76), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n460_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT10), .B(G99gat), .Z(new_n493_));
  INV_X1    g292(.A(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G85gat), .B(G92gat), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT9), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n495_), .B(new_n497_), .C1(KEYINPUT9), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n502_), .A2(KEYINPUT64), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT64), .B1(new_n502_), .B2(new_n503_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT66), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514_));
  INV_X1    g313(.A(G99gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n494_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT66), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n510_), .ZN(new_n518_));
  AND3_X1   g317(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT65), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n502_), .A2(new_n522_), .A3(new_n503_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n513_), .A2(new_n518_), .A3(new_n521_), .A4(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n496_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT67), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT8), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT8), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n496_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n511_), .A2(new_n512_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n506_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n528_), .B1(new_n524_), .B2(new_n496_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(new_n526_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n509_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT12), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT11), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n538_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(KEYINPUT11), .B2(new_n539_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT68), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n540_), .A2(new_n541_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n536_), .A2(new_n537_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n531_), .B1(new_n534_), .B2(new_n526_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n496_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n516_), .A2(new_n517_), .A3(new_n510_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n517_), .B1(new_n516_), .B2(new_n510_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n521_), .A2(new_n523_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n555_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT67), .B1(new_n560_), .B2(new_n528_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n508_), .B1(new_n554_), .B2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT12), .B1(new_n562_), .B2(new_n551_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n553_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n562_), .B2(new_n551_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n536_), .A2(new_n552_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n551_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n564_), .A2(new_n567_), .B1(new_n570_), .B2(new_n566_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT70), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT13), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT69), .B1(new_n571_), .B2(new_n576_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n537_), .B1(new_n536_), .B2(new_n552_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n562_), .A2(KEYINPUT12), .A3(new_n551_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n567_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n570_), .A2(new_n566_), .ZN(new_n584_));
  AND4_X1   g383(.A1(KEYINPUT69), .A2(new_n583_), .A3(new_n584_), .A4(new_n576_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n577_), .B(new_n579_), .C1(new_n580_), .C2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n578_), .A2(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n584_), .A3(new_n576_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT69), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n571_), .A2(KEYINPUT69), .A3(new_n576_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n587_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(new_n577_), .A3(new_n579_), .A4(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT72), .ZN(new_n599_));
  XOR2_X1   g398(.A(G134gat), .B(G162gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT36), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT34), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT35), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n536_), .A2(KEYINPUT71), .A3(new_n480_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT71), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n562_), .B2(new_n479_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n472_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n562_), .A2(new_n614_), .B1(new_n607_), .B2(new_n606_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n609_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n613_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n603_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n601_), .A2(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n620_), .A2(new_n622_), .A3(new_n616_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n597_), .B1(new_n619_), .B2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n602_), .B1(new_n620_), .B2(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n617_), .A2(new_n618_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n625_), .B(KEYINPUT37), .C1(new_n626_), .C2(new_n622_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n467_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n551_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631_));
  XOR2_X1   g430(.A(G127gat), .B(G155gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT16), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n630_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(KEYINPUT17), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n630_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT73), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n624_), .A2(new_n627_), .A3(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n596_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT74), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n492_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n644_), .A2(G1gat), .A3(new_n300_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT101), .Z(new_n647_));
  NOR2_X1   g446(.A1(new_n619_), .A2(new_n623_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n460_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n490_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n596_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT102), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n639_), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n300_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n647_), .B(new_n655_), .C1(KEYINPUT38), .C2(new_n645_), .ZN(G1324gat));
  NAND4_X1  g455(.A1(new_n492_), .A2(new_n463_), .A3(new_n428_), .A4(new_n643_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n654_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n463_), .B1(new_n658_), .B2(new_n428_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT40), .B(new_n657_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  INV_X1    g466(.A(new_n440_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G15gat), .B1(new_n654_), .B2(new_n668_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n669_), .A2(KEYINPUT41), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(KEYINPUT41), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n440_), .A2(new_n208_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n670_), .B(new_n671_), .C1(new_n644_), .C2(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(new_n362_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G22gat), .B1(new_n654_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n674_), .A2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n644_), .B2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(new_n640_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n648_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT104), .Z(new_n681_));
  INV_X1    g480(.A(new_n596_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n492_), .A2(new_n683_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n684_), .A2(G29gat), .A3(new_n300_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n624_), .A2(new_n627_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n436_), .B2(new_n459_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT43), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n689_), .B(new_n686_), .C1(new_n436_), .C2(new_n459_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n640_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n653_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT44), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n299_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n693_), .B2(new_n299_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n685_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  XOR2_X1   g497(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n684_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n434_), .A2(G36gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NOR4_X1   g502(.A1(new_n684_), .A2(G36gat), .A3(new_n434_), .A4(new_n699_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n693_), .A2(new_n428_), .ZN(new_n706_));
  INV_X1    g505(.A(G36gat), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT46), .B(new_n705_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n693_), .B2(new_n428_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n705_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(G1329gat));
  NOR3_X1   g512(.A1(new_n684_), .A2(G43gat), .A3(new_n668_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n693_), .A2(new_n258_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT47), .B(new_n715_), .C1(new_n716_), .C2(new_n212_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n212_), .B1(new_n693_), .B2(new_n258_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n714_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1330gat));
  NAND2_X1  g520(.A1(new_n693_), .A2(new_n362_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G50gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n674_), .A2(G50gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT106), .Z(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n684_), .B2(new_n725_), .ZN(G1331gat));
  INV_X1    g525(.A(new_n491_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n650_), .A2(new_n727_), .A3(new_n640_), .A4(new_n596_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n300_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n682_), .A2(new_n490_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n460_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n686_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n640_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n300_), .A2(G57gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1332gat));
  OAI21_X1  g534(.A(G64gat), .B1(new_n728_), .B2(new_n434_), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n434_), .A2(G64gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n733_), .B2(new_n739_), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n728_), .B2(new_n668_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n668_), .A2(G71gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n733_), .B2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n728_), .B2(new_n674_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n747_));
  OR2_X1    g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n747_), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n733_), .A2(G78gat), .A3(new_n674_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n731_), .A2(new_n681_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(G85gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n299_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n691_), .A2(new_n730_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n299_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n757_), .B2(new_n754_), .ZN(G1336gat));
  INV_X1    g557(.A(G92gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n759_), .A3(new_n428_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n756_), .A2(new_n428_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n759_), .ZN(G1337gat));
  AOI21_X1  g561(.A(new_n515_), .B1(new_n756_), .B2(new_n440_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n258_), .A2(new_n493_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n753_), .B2(new_n764_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g565(.A1(new_n753_), .A2(new_n494_), .A3(new_n362_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n691_), .A2(KEYINPUT110), .A3(new_n362_), .A4(new_n730_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(G106gat), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n688_), .A2(new_n690_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(new_n362_), .A3(new_n679_), .A4(new_n730_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n768_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  AND4_X1   g574(.A1(new_n768_), .A2(new_n774_), .A3(G106gat), .A4(new_n769_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n767_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n767_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  XOR2_X1   g580(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n642_), .B2(new_n727_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n596_), .A2(new_n641_), .A3(new_n491_), .A4(new_n782_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n787_));
  NAND2_X1  g586(.A1(new_n593_), .A2(new_n577_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n473_), .A2(new_n482_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n481_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n487_), .B(new_n789_), .C1(new_n790_), .C2(new_n482_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n488_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT55), .B(new_n567_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n583_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n569_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n566_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n564_), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n567_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n798_), .A2(new_n800_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n795_), .B(KEYINPUT56), .C1(new_n804_), .C2(new_n575_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n593_), .A2(new_n490_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n575_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n795_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n794_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n787_), .B1(new_n813_), .B2(new_n648_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n795_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n575_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n806_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n808_), .A2(KEYINPUT113), .A3(new_n809_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n793_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT57), .A3(new_n649_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n810_), .A2(new_n811_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n792_), .A2(new_n593_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT58), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n686_), .A3(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n814_), .A2(new_n822_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n639_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n786_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n258_), .A2(new_n299_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT59), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n812_), .A2(new_n819_), .A3(new_n818_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n648_), .B1(new_n838_), .B2(new_n793_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n732_), .B1(new_n827_), .B2(KEYINPUT58), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n839_), .A2(KEYINPUT57), .B1(new_n826_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n640_), .B1(new_n841_), .B2(new_n814_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n837_), .B1(new_n842_), .B2(new_n786_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT115), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n836_), .A2(new_n843_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n727_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n832_), .A2(new_n835_), .ZN(new_n850_));
  INV_X1    g649(.A(G113gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n490_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(G1340gat));
  OAI21_X1  g652(.A(G120gat), .B1(new_n844_), .B2(new_n682_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n596_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n850_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n854_), .A2(new_n859_), .ZN(G1341gat));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n836_), .A2(new_n846_), .A3(new_n843_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n846_), .B1(new_n836_), .B2(new_n843_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT116), .B(G127gat), .Z(new_n864_));
  NAND2_X1  g663(.A1(new_n639_), .A2(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n862_), .A2(new_n863_), .A3(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n832_), .A2(new_n679_), .A3(new_n835_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(G127gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n861_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n868_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT117), .B(new_n870_), .C1(new_n848_), .C2(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n848_), .B2(new_n732_), .ZN(new_n873_));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n850_), .A2(new_n874_), .A3(new_n648_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n668_), .A2(new_n362_), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n832_), .A2(new_n300_), .A3(new_n428_), .A4(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n490_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n596_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n640_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  AOI21_X1  g684(.A(G162gat), .B1(new_n878_), .B2(new_n648_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n686_), .A2(G162gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT118), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n878_), .B2(new_n888_), .ZN(G1347gat));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n830_), .A2(new_n679_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n786_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n434_), .A2(new_n299_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n440_), .A2(new_n894_), .A3(new_n674_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n651_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n890_), .B1(new_n898_), .B2(new_n230_), .ZN(new_n899_));
  OAI211_X1 g698(.A(KEYINPUT62), .B(G169gat), .C1(new_n897_), .C2(new_n651_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n370_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT119), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n899_), .A2(new_n904_), .A3(new_n900_), .A4(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1348gat));
  NOR2_X1   g705(.A1(new_n832_), .A2(new_n895_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(G176gat), .A3(new_n596_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT120), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n895_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G176gat), .B1(new_n910_), .B2(new_n596_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1349gat));
  NOR3_X1   g711(.A1(new_n897_), .A2(new_n235_), .A3(new_n831_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G183gat), .B1(new_n907_), .B2(new_n640_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n897_), .B2(new_n732_), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(KEYINPUT121), .Z(new_n917_));
  NAND3_X1  g716(.A1(new_n648_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT122), .Z(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n897_), .B2(new_n919_), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n832_), .A2(new_n877_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n921_), .A2(G197gat), .A3(new_n490_), .A4(new_n894_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n921_), .A2(new_n894_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n490_), .ZN(new_n926_));
  INV_X1    g725(.A(G197gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT124), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n926_), .A2(new_n930_), .A3(new_n927_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n924_), .B1(new_n929_), .B2(new_n931_), .ZN(G1352gat));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n682_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n925_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(G204gat), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n921_), .A2(new_n894_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n935_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT126), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  AND4_X1   g739(.A1(new_n933_), .A2(new_n936_), .A3(new_n937_), .A4(new_n940_), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n936_), .A2(new_n940_), .B1(new_n933_), .B2(new_n937_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1353gat));
  NOR2_X1   g742(.A1(new_n938_), .A2(new_n831_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  AND2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(new_n944_), .B2(new_n945_), .ZN(G1354gat));
  XOR2_X1   g747(.A(KEYINPUT127), .B(G218gat), .Z(new_n949_));
  NOR3_X1   g748(.A1(new_n938_), .A2(new_n732_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n925_), .A2(new_n648_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n949_), .ZN(G1355gat));
endmodule


