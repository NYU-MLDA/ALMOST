//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n213_), .B(new_n214_), .Z(new_n215_));
  XNOR2_X1  g014(.A(new_n208_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(new_n215_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n221_));
  INV_X1    g020(.A(new_n215_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n223_), .A3(new_n217_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G141gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G197gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n219_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n238_));
  OAI21_X1  g037(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n239_));
  OR3_X1    g038(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n235_), .A2(G183gat), .A3(G190gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n242_), .A2(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT24), .A3(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT26), .B(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n253_));
  INV_X1    g052(.A(G183gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(KEYINPUT25), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT25), .B(G183gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n252_), .B(new_n255_), .C1(new_n256_), .C2(new_n253_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n248_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n246_), .A2(new_n247_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n241_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT81), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT30), .Z(new_n263_));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT84), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n265_), .B(new_n269_), .Z(new_n270_));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(G15gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G71gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G99gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(KEYINPUT82), .B(G43gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT31), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n270_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT85), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(KEYINPUT2), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT86), .B1(new_n289_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n287_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT86), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n286_), .B1(new_n297_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n285_), .B1(new_n283_), .B2(KEYINPUT1), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(KEYINPUT1), .B2(new_n285_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n291_), .A2(new_n292_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n306_), .A2(new_n299_), .A3(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT28), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G211gat), .B(G218gat), .Z(new_n314_));
  INV_X1    g113(.A(KEYINPUT21), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT21), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n314_), .A3(KEYINPUT21), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT88), .ZN(new_n323_));
  AND2_X1   g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n324_), .A2(new_n323_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n325_), .B(new_n329_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n328_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n313_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G22gat), .B(G50gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n330_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n328_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n339_), .A2(new_n332_), .A3(new_n312_), .A4(new_n331_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n335_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n256_), .A2(new_n252_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT89), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT90), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n250_), .B(new_n238_), .C1(new_n349_), .C2(G176gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n322_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT91), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n322_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n262_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n353_), .A2(KEYINPUT20), .A3(new_n355_), .A4(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n347_), .A2(new_n350_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n354_), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT20), .B(new_n361_), .C1(new_n262_), .C2(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n357_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT93), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n364_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n359_), .B2(new_n363_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n269_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n309_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n268_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT4), .B(new_n379_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n385_), .A2(new_n383_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n269_), .B(new_n387_), .C1(new_n304_), .C2(new_n308_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT94), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n384_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n372_), .A2(new_n373_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n383_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n382_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(new_n393_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n394_), .B(new_n377_), .C1(new_n389_), .C2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT95), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT33), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(KEYINPUT95), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n392_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n394_), .B1(new_n389_), .B2(new_n395_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n378_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n396_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n362_), .A2(new_n357_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n322_), .A2(new_n346_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(new_n350_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n358_), .B1(new_n355_), .B2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n412_));
  MUX2_X1   g211(.A(new_n411_), .B(new_n364_), .S(new_n412_), .Z(new_n413_));
  AOI22_X1  g212(.A1(new_n401_), .A2(new_n402_), .B1(new_n405_), .B2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n392_), .A2(new_n398_), .A3(KEYINPUT96), .A4(new_n400_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n344_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n405_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n372_), .A2(KEYINPUT27), .A3(new_n373_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT98), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n364_), .B2(new_n371_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n359_), .A2(new_n363_), .A3(KEYINPUT98), .A4(new_n370_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n421_), .B(new_n422_), .C1(new_n370_), .C2(new_n411_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n423_), .B2(KEYINPUT27), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n282_), .B1(new_n416_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n344_), .A2(new_n424_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n417_), .A3(new_n281_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n233_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G57gat), .B(G64gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT11), .ZN(new_n431_));
  XOR2_X1   g230(.A(G71gat), .B(G78gat), .Z(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n431_), .A2(new_n432_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n430_), .A2(KEYINPUT11), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n433_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438_));
  INV_X1    g237(.A(G85gat), .ZN(new_n439_));
  INV_X1    g238(.A(G92gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT64), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT64), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G92gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n439_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n444_), .B2(KEYINPUT9), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT9), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT64), .B(G92gat), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT65), .B(new_n446_), .C1(new_n447_), .C2(new_n439_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G85gat), .B(G92gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(KEYINPUT9), .B2(new_n440_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n445_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n445_), .A2(KEYINPUT66), .A3(new_n448_), .A4(new_n450_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT10), .B(G99gat), .Z(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT6), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n453_), .A2(new_n454_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  INV_X1    g265(.A(new_n449_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT67), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT7), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(new_n470_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n459_), .A2(new_n461_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n466_), .B(new_n467_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n471_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT67), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n470_), .B1(new_n469_), .B2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n459_), .A2(new_n461_), .A3(KEYINPUT68), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT68), .B1(new_n459_), .B2(new_n461_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n467_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n476_), .B1(new_n487_), .B2(KEYINPUT8), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT12), .B(new_n437_), .C1(new_n465_), .C2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT71), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n437_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n473_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT8), .B1(new_n493_), .B2(new_n449_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n475_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n453_), .A2(new_n454_), .A3(new_n464_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT72), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n497_), .B2(KEYINPUT12), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n463_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n454_), .A2(new_n503_), .B1(new_n494_), .B2(new_n475_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT72), .B(new_n502_), .C1(new_n504_), .C2(new_n492_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(G230gat), .A2(G233gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n504_), .B2(new_n492_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n499_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n497_), .A2(KEYINPUT70), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n504_), .B2(new_n492_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n495_), .A2(new_n496_), .A3(new_n492_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT69), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n504_), .A2(KEYINPUT69), .A3(new_n492_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n510_), .A2(new_n512_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n507_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G120gat), .B(G148gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT5), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G176gat), .B(G204gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n509_), .A2(new_n518_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n527_), .B(KEYINPUT13), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT73), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n495_), .A2(new_n496_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n221_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n504_), .A2(new_n206_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT75), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n537_), .A2(new_n538_), .A3(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n537_), .A2(new_n538_), .A3(new_n547_), .A4(new_n543_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(KEYINPUT74), .A3(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G134gat), .B(G162gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n549_), .B(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n546_), .A2(new_n548_), .ZN(new_n556_));
  OR3_X1    g355(.A1(new_n556_), .A2(new_n553_), .A3(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT76), .A3(KEYINPUT37), .ZN(new_n559_));
  OR2_X1    g358(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n560_));
  NAND2_X1  g359(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n555_), .A2(new_n557_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n215_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n492_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n571_), .B2(KEYINPUT17), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(KEYINPUT17), .B2(new_n568_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n575_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AND4_X1   g378(.A1(new_n429_), .A2(new_n535_), .A3(new_n564_), .A4(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n210_), .A3(new_n405_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n580_), .A2(KEYINPUT99), .A3(new_n210_), .A4(new_n405_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(KEYINPUT38), .A3(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n558_), .B(KEYINPUT101), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n535_), .A2(new_n232_), .A3(new_n579_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n587_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n417_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n583_), .A2(new_n584_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT102), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n597_), .B(KEYINPUT38), .C1(new_n583_), .C2(new_n584_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n585_), .B(new_n593_), .C1(new_n596_), .C2(new_n598_), .ZN(G1324gat));
  NAND3_X1  g398(.A1(new_n580_), .A2(new_n211_), .A3(new_n424_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n424_), .B(new_n587_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n211_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n600_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n606_), .B(new_n608_), .ZN(G1325gat));
  NAND3_X1  g408(.A1(new_n580_), .A2(new_n272_), .A3(new_n281_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n592_), .A2(new_n282_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n611_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(new_n611_), .B2(G15gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n612_), .B2(new_n613_), .ZN(G1326gat));
  INV_X1    g413(.A(G22gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n580_), .A2(new_n615_), .A3(new_n344_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G22gat), .B1(new_n592_), .B2(new_n343_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(KEYINPUT42), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(KEYINPUT42), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n616_), .B1(new_n618_), .B2(new_n619_), .ZN(G1327gat));
  NAND4_X1  g419(.A1(new_n533_), .A2(new_n531_), .A3(new_n232_), .A4(new_n578_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT105), .Z(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(KEYINPUT106), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n564_), .B(new_n624_), .C1(new_n426_), .C2(new_n428_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n401_), .A2(new_n402_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n413_), .A2(new_n405_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n415_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n425_), .B1(new_n629_), .B2(new_n343_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n428_), .B1(new_n630_), .B2(new_n281_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n626_), .B1(new_n631_), .B2(new_n563_), .ZN(new_n632_));
  OAI211_X1 g431(.A(KEYINPUT44), .B(new_n622_), .C1(new_n625_), .C2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n624_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(new_n563_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n564_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(new_n626_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT44), .B1(new_n638_), .B2(new_n622_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n634_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n405_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G29gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n578_), .A2(new_n558_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n534_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n429_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n417_), .A2(G29gat), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT107), .Z(new_n648_));
  OAI21_X1  g447(.A(new_n642_), .B1(new_n646_), .B2(new_n648_), .ZN(G1328gat));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  INV_X1    g449(.A(G36gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n640_), .B2(new_n424_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n651_), .A3(new_n424_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT45), .Z(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n653_), .B(KEYINPUT45), .ZN(new_n656_));
  INV_X1    g455(.A(new_n424_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n634_), .A2(new_n639_), .A3(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n656_), .B(KEYINPUT46), .C1(new_n658_), .C2(new_n651_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(G1329gat));
  AND2_X1   g459(.A1(new_n281_), .A2(G43gat), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n640_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT108), .B(G43gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n646_), .B2(new_n282_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT47), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT47), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(new_n667_), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1330gat));
  AOI21_X1  g468(.A(G50gat), .B1(new_n645_), .B2(new_n344_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n344_), .A2(G50gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n640_), .B2(new_n671_), .ZN(G1331gat));
  NOR2_X1   g471(.A1(new_n578_), .A2(new_n232_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n587_), .A2(new_n534_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n405_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G57gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n232_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n535_), .A2(new_n563_), .A3(new_n578_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n417_), .A2(G57gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g483(.A(G64gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n674_), .B2(new_n424_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT48), .Z(new_n687_));
  INV_X1    g486(.A(new_n681_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n685_), .A3(new_n424_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1333gat));
  AOI21_X1  g489(.A(new_n274_), .B1(new_n674_), .B2(new_n281_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n281_), .A2(new_n274_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n681_), .B2(new_n694_), .ZN(G1334gat));
  INV_X1    g494(.A(G78gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n674_), .B2(new_n344_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT50), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n688_), .A2(new_n696_), .A3(new_n344_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1335gat));
  NOR3_X1   g499(.A1(new_n535_), .A2(new_n232_), .A3(new_n579_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n638_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n405_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G85gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n535_), .A2(new_n643_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n679_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n405_), .A2(new_n439_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(new_n440_), .B1(new_n706_), .B2(new_n657_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n657_), .A2(new_n447_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n711_), .A2(new_n712_), .B1(new_n702_), .B2(new_n713_), .ZN(G1337gat));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(KEYINPUT51), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n638_), .A2(new_n281_), .A3(new_n701_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G99gat), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n679_), .A2(new_n281_), .A3(new_n455_), .A4(new_n705_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n715_), .A2(KEYINPUT51), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n638_), .A2(new_n344_), .A3(new_n701_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G106gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G106gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n344_), .A2(new_n456_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n725_), .A2(new_n726_), .B1(new_n706_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT53), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730_));
  OAI221_X1 g529(.A(new_n730_), .B1(new_n706_), .B2(new_n727_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1339gat));
  INV_X1    g531(.A(G113gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n216_), .A2(new_n217_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n220_), .A2(new_n223_), .A3(new_n218_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n229_), .A3(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n526_), .A2(new_n231_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n499_), .A2(new_n506_), .A3(new_n513_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n507_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n509_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n499_), .A2(new_n506_), .A3(KEYINPUT55), .A4(new_n508_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n743_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT56), .B1(new_n743_), .B2(new_n523_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n737_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT58), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT58), .B(new_n737_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n563_), .A3(new_n749_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n526_), .A2(KEYINPUT114), .A3(new_n232_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT114), .B1(new_n526_), .B2(new_n232_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n527_), .A2(new_n231_), .A3(new_n736_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n558_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n750_), .B1(KEYINPUT57), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(KEYINPUT57), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n579_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n564_), .A2(new_n532_), .A3(new_n673_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n427_), .A2(new_n405_), .A3(new_n281_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n733_), .B1(new_n767_), .B2(new_n233_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(KEYINPUT59), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n563_), .A2(new_n749_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n743_), .A2(new_n523_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n743_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT58), .B1(new_n778_), .B2(new_n737_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n773_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n754_), .A2(new_n755_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n558_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT57), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n772_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n750_), .B(KEYINPUT116), .C1(KEYINPUT57), .C2(new_n756_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n759_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n763_), .B1(new_n786_), .B2(new_n578_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n765_), .A2(KEYINPUT59), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n771_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n232_), .A2(G113gat), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT117), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n769_), .A2(new_n770_), .B1(new_n792_), .B2(new_n794_), .ZN(G1340gat));
  XNOR2_X1  g594(.A(KEYINPUT118), .B(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n791_), .B2(new_n535_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT60), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n534_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT119), .B1(new_n796_), .B2(new_n798_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n797_), .B1(new_n767_), .B2(new_n803_), .ZN(G1341gat));
  OAI21_X1  g603(.A(G127gat), .B1(new_n791_), .B2(new_n578_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n578_), .A2(G127gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n767_), .B2(new_n806_), .ZN(G1342gat));
  OAI21_X1  g606(.A(G134gat), .B1(new_n791_), .B2(new_n564_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n586_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(G134gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n767_), .B2(new_n810_), .ZN(G1343gat));
  NOR3_X1   g610(.A1(new_n281_), .A2(new_n417_), .A3(new_n343_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n764_), .A2(new_n657_), .A3(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n233_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(new_n291_), .ZN(G1344gat));
  NOR2_X1   g614(.A1(new_n813_), .A2(new_n535_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT120), .B(G148gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1345gat));
  NOR2_X1   g617(.A1(new_n813_), .A2(new_n578_), .ZN(new_n819_));
  XOR2_X1   g618(.A(KEYINPUT61), .B(G155gat), .Z(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  OAI21_X1  g620(.A(G162gat), .B1(new_n813_), .B2(new_n564_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n809_), .A2(G162gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n813_), .B2(new_n823_), .ZN(G1347gat));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n282_), .A2(new_n657_), .A3(new_n344_), .A4(new_n405_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n759_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n757_), .B2(new_n772_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n579_), .B1(new_n828_), .B2(new_n785_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n232_), .B(new_n826_), .C1(new_n829_), .C2(new_n763_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G169gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n825_), .B1(new_n831_), .B2(KEYINPUT62), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(KEYINPUT62), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n830_), .A2(KEYINPUT121), .A3(new_n834_), .A4(G169gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n837_));
  INV_X1    g636(.A(new_n826_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n787_), .B2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT122), .B(new_n826_), .C1(new_n829_), .C2(new_n763_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n349_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n232_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(new_n843_), .ZN(G1348gat));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  AOI21_X1  g644(.A(G176gat), .B1(new_n841_), .B2(new_n534_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n764_), .A2(G176gat), .A3(new_n534_), .A4(new_n826_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n535_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n847_), .B(KEYINPUT123), .C1(new_n850_), .C2(G176gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1349gat));
  NOR2_X1   g651(.A1(new_n760_), .A2(new_n763_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n853_), .A2(new_n578_), .A3(new_n838_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n854_), .A2(KEYINPUT124), .ZN(new_n855_));
  AOI21_X1  g654(.A(G183gat), .B1(new_n854_), .B2(KEYINPUT124), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n578_), .A2(new_n256_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n855_), .A2(new_n856_), .B1(new_n841_), .B2(new_n857_), .ZN(G1350gat));
  NAND3_X1  g657(.A1(new_n841_), .A2(new_n252_), .A3(new_n586_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n564_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n860_));
  INV_X1    g659(.A(G190gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1351gat));
  OR3_X1    g661(.A1(new_n281_), .A2(new_n657_), .A3(new_n418_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n853_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n232_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n534_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g667(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n578_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n864_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n873_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n870_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n872_), .A2(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n873_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n869_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1354gat));
  NOR2_X1   g679(.A1(new_n809_), .A2(G218gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n864_), .A2(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n853_), .A2(new_n564_), .A3(new_n863_), .ZN(new_n883_));
  INV_X1    g682(.A(G218gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


