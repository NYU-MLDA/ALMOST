//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT91), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(G197gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT91), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(new_n205_), .A3(G197gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT21), .ZN(new_n212_));
  XOR2_X1   g011(.A(G211gat), .B(G218gat), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n206_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(KEYINPUT21), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n213_), .A2(KEYINPUT21), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n212_), .A2(new_n215_), .B1(new_n211_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT79), .B(G183gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT25), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(KEYINPUT25), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT81), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n219_), .A2(new_n229_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT23), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT82), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n233_), .B(new_n236_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n231_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G169gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT84), .ZN(new_n245_));
  AOI21_X1  g044(.A(G176gat), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT83), .B(G169gat), .Z(new_n247_));
  OAI221_X1 g046(.A(new_n246_), .B1(new_n245_), .B2(new_n244_), .C1(new_n247_), .C2(new_n243_), .ZN(new_n248_));
  INV_X1    g047(.A(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n218_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n233_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n238_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n217_), .B1(new_n242_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n233_), .A2(new_n236_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT95), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n237_), .A2(KEYINPUT24), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT94), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n234_), .B1(new_n258_), .B2(KEYINPUT94), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT25), .B(G183gat), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n259_), .A2(new_n260_), .B1(new_n226_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n233_), .A2(KEYINPUT95), .A3(new_n236_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n233_), .B1(G183gat), .B2(G190gat), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT22), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n244_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n265_), .B(new_n252_), .C1(G176gat), .C2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n212_), .A2(new_n215_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n216_), .A2(new_n211_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT20), .B1(new_n270_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n204_), .B1(new_n254_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n276_), .B1(new_n270_), .B2(new_n273_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n242_), .A2(new_n253_), .A3(new_n217_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n203_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT18), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(new_n278_), .A3(new_n204_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n254_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT99), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n270_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n264_), .A2(KEYINPUT99), .A3(new_n269_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n217_), .A3(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n288_), .B1(new_n295_), .B2(new_n203_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n286_), .B(KEYINPUT27), .C1(new_n296_), .C2(new_n285_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n280_), .A2(new_n285_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n284_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G127gat), .B(G134gat), .Z(new_n305_));
  XOR2_X1   g104(.A(G113gat), .B(G120gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT96), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n316_));
  OR2_X1    g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(KEYINPUT3), .ZN(new_n318_));
  NOR3_X1   g117(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT89), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n315_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(G155gat), .A3(G162gat), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT88), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(KEYINPUT1), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n329_), .A2(new_n327_), .A3(new_n322_), .A4(KEYINPUT88), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n328_), .A2(new_n330_), .A3(new_n317_), .A4(new_n310_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n308_), .B(new_n309_), .C1(new_n325_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n324_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n318_), .A2(new_n320_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n315_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n307_), .A3(new_n331_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n333_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n304_), .B(new_n335_), .C1(new_n340_), .C2(new_n334_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n307_), .B1(new_n338_), .B2(new_n331_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n303_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT100), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT100), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n341_), .A2(new_n351_), .A3(new_n345_), .A4(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n341_), .A2(new_n348_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n345_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n302_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G78gat), .B(G106gat), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n331_), .B(new_n360_), .C1(new_n321_), .C2(new_n324_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT28), .A2(G22gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G50gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(KEYINPUT28), .A2(G22gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(G50gat), .B1(new_n368_), .B2(new_n363_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n362_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n367_), .A2(new_n369_), .A3(new_n362_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n361_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n370_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n373_), .A2(new_n338_), .A3(new_n360_), .A4(new_n331_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n360_), .B1(new_n338_), .B2(new_n331_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n217_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT29), .B1(new_n325_), .B2(new_n332_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n273_), .A3(new_n377_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT93), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n375_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n376_), .A2(new_n380_), .A3(new_n387_), .A4(new_n382_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n359_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G43gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT86), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n242_), .A2(new_n253_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n253_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n240_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(G71gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G99gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n395_), .A2(new_n398_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT87), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n395_), .A2(new_n398_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n406_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n307_), .B(KEYINPUT31), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT87), .B(new_n417_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n384_), .A2(new_n388_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n385_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n358_), .A3(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n391_), .A2(new_n419_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n419_), .B1(new_n391_), .B2(new_n423_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n357_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n295_), .A2(new_n203_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n285_), .A2(KEYINPUT32), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n287_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT97), .B1(new_n275_), .B2(new_n279_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n432_));
  OAI22_X1  g231(.A1(new_n429_), .A2(new_n430_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n356_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n299_), .A2(new_n300_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n340_), .A2(new_n334_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n335_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n303_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n346_), .A2(new_n347_), .A3(new_n303_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n345_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n442_));
  AOI211_X1 g241(.A(KEYINPUT33), .B(new_n345_), .C1(new_n341_), .C2(new_n348_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n435_), .B(new_n440_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n444_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n391_), .A2(new_n423_), .B1(new_n418_), .B2(new_n416_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n426_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G230gat), .A2(G233gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n449_), .B(KEYINPUT64), .Z(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT9), .A3(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(KEYINPUT9), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n454_), .A2(new_n458_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT7), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(new_n402_), .A3(new_n456_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT65), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n464_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n466_), .A2(new_n454_), .A3(new_n467_), .A4(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n459_), .A2(new_n460_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n472_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n463_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G57gat), .B(G64gat), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n480_));
  XOR2_X1   g279(.A(G71gat), .B(G78gat), .Z(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n477_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n484_), .B(new_n463_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(KEYINPUT12), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n477_), .A2(new_n489_), .A3(new_n485_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n451_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n450_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G120gat), .B(G148gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT5), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G176gat), .B(G204gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  NOR3_X1   g295(.A1(new_n491_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT13), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(KEYINPUT13), .A3(new_n499_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G29gat), .B(G36gat), .Z(new_n505_));
  XOR2_X1   g304(.A(G43gat), .B(G50gat), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G29gat), .B(G36gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G43gat), .B(G50gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n507_), .A2(KEYINPUT15), .A3(new_n510_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516_));
  INV_X1    g315(.A(G1gat), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G8gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n511_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n522_), .B(new_n524_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G113gat), .B(G141gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT78), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G169gat), .B(G197gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n504_), .A2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n448_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT17), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n484_), .B(new_n522_), .ZN(new_n550_));
  AND2_X1   g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n546_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n463_), .B(new_n511_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT34), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT67), .ZN(new_n565_));
  INV_X1    g364(.A(new_n463_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT6), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n467_), .ZN(new_n571_));
  NOR4_X1   g370(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n469_), .B1(new_n468_), .B2(new_n464_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n474_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT8), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n566_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n513_), .A2(new_n514_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n565_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n477_), .A2(new_n515_), .A3(KEYINPUT67), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n564_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT68), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n560_), .A2(new_n563_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n578_), .A2(new_n565_), .A3(new_n579_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT67), .B1(new_n477_), .B2(new_n515_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT68), .ZN(new_n589_));
  INV_X1    g388(.A(new_n583_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n583_), .B(KEYINPUT70), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n585_), .B(new_n593_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n582_), .A2(KEYINPUT71), .A3(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT69), .ZN(new_n600_));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(KEYINPUT36), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n592_), .A2(new_n598_), .A3(new_n603_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n584_), .A2(new_n591_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n602_), .B(KEYINPUT36), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n541_), .A2(new_n559_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n356_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT102), .Z(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT72), .B1(new_n605_), .B2(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n592_), .A2(new_n598_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT72), .ZN(new_n614_));
  INV_X1    g413(.A(new_n606_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n616_), .A3(new_n604_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT37), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n617_), .B2(KEYINPUT37), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n607_), .A2(KEYINPUT37), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n554_), .A2(KEYINPUT77), .A3(new_n557_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT77), .B1(new_n554_), .B2(new_n557_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n541_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT101), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n609_), .A2(G1gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(KEYINPUT38), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n611_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT38), .B1(new_n629_), .B2(new_n630_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT103), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n629_), .A2(new_n518_), .A3(new_n302_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n302_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G8gat), .B1(new_n608_), .B2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n636_), .B(new_n640_), .C1(new_n638_), .C2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g442(.A(G15gat), .B1(new_n608_), .B2(new_n419_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT41), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n628_), .A2(G15gat), .A3(new_n419_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1326gat));
  NAND2_X1  g446(.A1(new_n391_), .A2(new_n423_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G22gat), .B1(new_n608_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT42), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n648_), .A2(G22gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n628_), .B2(new_n651_), .ZN(G1327gat));
  NOR2_X1   g451(.A1(new_n625_), .A2(new_n607_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n541_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G29gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n356_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n606_), .B1(new_n592_), .B2(new_n598_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n604_), .B1(new_n659_), .B2(new_n614_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n605_), .A2(KEYINPUT72), .A3(new_n606_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT37), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n621_), .B1(new_n662_), .B2(KEYINPUT73), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT37), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n448_), .A3(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT105), .B1(new_n665_), .B2(KEYINPUT43), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(KEYINPUT43), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n540_), .A2(new_n626_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n658_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(KEYINPUT43), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n668_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n665_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n670_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(KEYINPUT44), .A3(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n671_), .A2(new_n356_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT106), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n671_), .A2(new_n679_), .A3(new_n682_), .A4(new_n356_), .ZN(new_n683_));
  AND4_X1   g482(.A1(KEYINPUT107), .A2(new_n681_), .A3(G29gat), .A4(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n656_), .B1(new_n680_), .B2(KEYINPUT106), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT107), .B1(new_n685_), .B2(new_n683_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n657_), .B1(new_n684_), .B2(new_n686_), .ZN(G1328gat));
  NAND2_X1  g486(.A1(new_n671_), .A2(new_n679_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G36gat), .B1(new_n688_), .B2(new_n637_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n654_), .A2(G36gat), .A3(new_n637_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT45), .Z(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n689_), .A2(KEYINPUT46), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1329gat));
  INV_X1    g495(.A(new_n419_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n671_), .A2(new_n679_), .A3(G43gat), .A4(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G43gat), .B1(new_n655_), .B2(new_n697_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT108), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(KEYINPUT108), .B2(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT47), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n701_), .B(new_n704_), .C1(KEYINPUT108), .C2(new_n698_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1330gat));
  OAI21_X1  g505(.A(G50gat), .B1(new_n688_), .B2(new_n648_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n648_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n365_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT109), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n654_), .B2(new_n710_), .ZN(G1331gat));
  NOR3_X1   g510(.A1(new_n623_), .A2(new_n624_), .A3(new_n538_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n448_), .A2(new_n607_), .A3(new_n504_), .A4(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n609_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n538_), .B1(new_n426_), .B2(new_n447_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT110), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n627_), .A3(new_n504_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n609_), .A2(G57gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n713_), .B2(new_n637_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT48), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n637_), .A2(G64gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n717_), .B2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n713_), .B2(new_n419_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n697_), .A2(new_n400_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n717_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n713_), .B2(new_n648_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n648_), .A2(G78gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n717_), .B2(new_n730_), .ZN(G1335gat));
  INV_X1    g530(.A(new_n607_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n716_), .A2(new_n626_), .A3(new_n732_), .A4(new_n504_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n356_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n504_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(new_n625_), .A3(new_n538_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n677_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n609_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1336gat));
  AOI21_X1  g541(.A(G92gat), .B1(new_n735_), .B2(new_n302_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n302_), .A2(G92gat), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT112), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n743_), .B1(new_n744_), .B2(new_n746_), .ZN(G1337gat));
  AOI21_X1  g546(.A(new_n402_), .B1(new_n744_), .B2(new_n697_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n697_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n735_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1338gat));
  XNOR2_X1  g551(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n677_), .A2(new_n708_), .A3(new_n739_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G106gat), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT52), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n735_), .A2(new_n456_), .A3(new_n708_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n754_), .B2(G106gat), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n757_), .B(new_n753_), .C1(new_n759_), .C2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n758_), .A2(new_n763_), .ZN(G1339gat));
  NAND2_X1  g563(.A1(new_n738_), .A2(new_n712_), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT54), .B(new_n765_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n662_), .A2(KEYINPUT73), .ZN(new_n768_));
  INV_X1    g567(.A(new_n621_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n664_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n765_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n766_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n498_), .A2(new_n538_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n488_), .A2(new_n451_), .A3(new_n490_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n491_), .B1(KEYINPUT55), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n488_), .A2(new_n490_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(KEYINPUT55), .A3(new_n450_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n496_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n775_), .A2(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n450_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n778_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n496_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n774_), .B1(new_n782_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n523_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n528_), .A2(new_n526_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n535_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n792_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n536_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n499_), .B2(new_n498_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n607_), .B1(new_n788_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT57), .B(new_n607_), .C1(new_n788_), .C2(new_n796_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n782_), .A2(KEYINPUT115), .A3(new_n787_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n795_), .A2(new_n497_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n782_), .B2(KEYINPUT115), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n802_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n782_), .A2(new_n787_), .A3(KEYINPUT115), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n496_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n807_), .A2(new_n810_), .A3(KEYINPUT58), .A4(new_n804_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n663_), .A2(new_n664_), .A3(new_n806_), .A4(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n559_), .B1(new_n801_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT116), .B1(new_n773_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n622_), .B2(new_n765_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n770_), .A2(new_n767_), .A3(new_n771_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n806_), .A2(new_n811_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n770_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n799_), .A2(new_n800_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n558_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n609_), .A2(new_n302_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n824_), .A2(new_n425_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n814_), .A2(new_n823_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT117), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n814_), .A2(new_n823_), .A3(new_n828_), .A4(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n538_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G113gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(KEYINPUT118), .A3(new_n831_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n825_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n626_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n817_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n836_), .B1(new_n837_), .B2(new_n842_), .ZN(new_n843_));
  AOI211_X1 g642(.A(KEYINPUT119), .B(new_n841_), .C1(new_n826_), .C2(KEYINPUT59), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n538_), .A2(G113gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT120), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n834_), .A2(new_n835_), .B1(new_n845_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  AOI21_X1  g648(.A(G120gat), .B1(new_n504_), .B2(new_n849_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT121), .Z(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n849_), .B2(G120gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n827_), .A2(new_n829_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT122), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n837_), .A2(new_n842_), .A3(new_n504_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G120gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n827_), .A2(new_n858_), .A3(new_n625_), .A4(new_n829_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n843_), .A2(new_n844_), .A3(new_n558_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n858_), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n827_), .A2(new_n862_), .A3(new_n732_), .A4(new_n829_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n843_), .A2(new_n844_), .A3(new_n770_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1343gat));
  AND2_X1   g664(.A1(new_n814_), .A2(new_n823_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n424_), .A3(new_n824_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n539_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT123), .B(G141gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1344gat));
  AND2_X1   g669(.A1(new_n866_), .A2(new_n424_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n504_), .A3(new_n824_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n867_), .A2(new_n626_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n867_), .B2(new_n770_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n607_), .A2(G162gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n867_), .B2(new_n878_), .ZN(G1347gat));
  NAND2_X1  g678(.A1(new_n817_), .A2(new_n840_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n637_), .A2(new_n356_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n697_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n708_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n266_), .B1(new_n885_), .B2(new_n538_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n538_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n887_), .B(new_n888_), .C1(new_n268_), .C2(new_n889_), .ZN(G1348gat));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n880_), .A2(new_n504_), .A3(new_n883_), .ZN(new_n892_));
  INV_X1    g691(.A(G176gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n892_), .A2(new_n891_), .A3(new_n893_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n866_), .A2(new_n648_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n881_), .A2(G176gat), .A3(new_n504_), .A4(new_n697_), .ZN(new_n897_));
  OAI22_X1  g696(.A1(new_n894_), .A2(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1349gat));
  NOR3_X1   g699(.A1(new_n884_), .A2(new_n558_), .A3(new_n261_), .ZN(new_n901_));
  OR3_X1    g700(.A1(new_n896_), .A2(new_n626_), .A3(new_n882_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n218_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n884_), .B2(new_n770_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n732_), .A2(new_n226_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n884_), .B2(new_n905_), .ZN(G1351gat));
  NAND3_X1  g705(.A1(new_n871_), .A2(new_n538_), .A3(new_n881_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT126), .B(G197gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1352gat));
  NAND3_X1  g708(.A1(new_n866_), .A2(new_n424_), .A3(new_n881_), .ZN(new_n910_));
  AND2_X1   g709(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n738_), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1353gat));
  XOR2_X1   g713(.A(KEYINPUT63), .B(G211gat), .Z(new_n915_));
  NAND4_X1  g714(.A1(new_n871_), .A2(new_n559_), .A3(new_n881_), .A4(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n910_), .B2(new_n558_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1354gat));
  OAI21_X1  g718(.A(G218gat), .B1(new_n910_), .B2(new_n770_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n607_), .A2(G218gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n910_), .B2(new_n921_), .ZN(G1355gat));
endmodule


