//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(new_n207_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G85gat), .B(G92gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n206_), .A2(new_n207_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n209_), .A2(new_n210_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT66), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n208_), .A2(new_n211_), .A3(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(KEYINPUT65), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT65), .B(KEYINPUT7), .Z(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(new_n229_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n226_), .A2(new_n228_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n223_), .B1(new_n234_), .B2(new_n220_), .ZN(new_n235_));
  AOI211_X1 g034(.A(KEYINPUT8), .B(new_n219_), .C1(new_n233_), .C2(new_n212_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n222_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G78gat), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G64gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(KEYINPUT11), .A3(new_n240_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n242_), .B(new_n243_), .C1(KEYINPUT11), .C2(new_n240_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n237_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n237_), .A2(new_n246_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(KEYINPUT68), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G230gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n237_), .A2(new_n252_), .A3(new_n246_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT5), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G176gat), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n244_), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT70), .B1(new_n248_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  AOI211_X1 g064(.A(new_n265_), .B(new_n262_), .C1(new_n237_), .C2(new_n246_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n261_), .B(new_n247_), .C1(new_n264_), .C2(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n254_), .B(new_n260_), .C1(new_n267_), .C2(new_n251_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT71), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n248_), .A2(new_n263_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n265_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n248_), .A2(KEYINPUT70), .A3(new_n263_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(new_n250_), .A3(new_n261_), .A4(new_n247_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n254_), .A4(new_n260_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n254_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n259_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT13), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT13), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n282_), .A3(new_n279_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT72), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(KEYINPUT72), .A3(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G29gat), .B(G36gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G43gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G50gat), .ZN(new_n292_));
  INV_X1    g091(.A(G43gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n290_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G50gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G22gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n301_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G8gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n297_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT77), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n297_), .A2(new_n307_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G229gat), .A2(G233gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT15), .B1(new_n292_), .B2(new_n296_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n292_), .A2(new_n296_), .A3(KEYINPUT15), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n307_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n309_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n312_), .B(KEYINPUT78), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n311_), .A2(new_n312_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G113gat), .B(G141gat), .ZN(new_n321_));
  INV_X1    g120(.A(G169gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G197gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  OAI221_X1 g126(.A(new_n327_), .B1(new_n318_), .B2(new_n319_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n287_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(KEYINPUT108), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n337_));
  XOR2_X1   g136(.A(G211gat), .B(G218gat), .Z(new_n338_));
  OR2_X1    g137(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n324_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n258_), .A2(G197gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(KEYINPUT21), .B(new_n338_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT95), .ZN(new_n344_));
  AND2_X1   g143(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(G197gat), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(G197gat), .B2(new_n258_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(KEYINPUT21), .A4(new_n338_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n324_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT93), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT21), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(G197gat), .B2(G204gat), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n347_), .B(new_n354_), .C1(G197gat), .C2(new_n258_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n338_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT94), .B1(new_n358_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(G197gat), .B1(new_n339_), .B2(new_n340_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT21), .B1(new_n324_), .B2(new_n258_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT93), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT92), .B(G204gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n342_), .B1(new_n368_), .B2(G197gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n338_), .B1(new_n369_), .B2(new_n354_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT94), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n351_), .B1(new_n362_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT23), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(G183gat), .A3(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT98), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n380_), .B(new_n382_), .C1(G176gat), .C2(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n388_), .B2(new_n381_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT26), .B(G190gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT25), .B(G183gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n374_), .A2(new_n393_), .A3(KEYINPUT23), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n375_), .A2(new_n377_), .A3(KEYINPUT82), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n389_), .A2(new_n392_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT107), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n385_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n397_), .B1(new_n385_), .B2(new_n396_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n337_), .B1(new_n373_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G190gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT79), .B1(new_n403_), .B2(KEYINPUT26), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(new_n391_), .C1(new_n390_), .C2(KEYINPUT79), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(new_n378_), .A3(new_n389_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n322_), .A2(KEYINPUT22), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT22), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G169gat), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT80), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT80), .B1(new_n409_), .B2(G169gat), .ZN(new_n412_));
  INV_X1    g211(.A(G176gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n407_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(G176gat), .B1(new_n408_), .B2(KEYINPUT80), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(KEYINPUT81), .C1(KEYINPUT80), .C2(new_n383_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n395_), .A2(new_n379_), .A3(new_n394_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n381_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n406_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT83), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(new_n406_), .C1(new_n418_), .C2(new_n420_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n344_), .A2(new_n350_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n367_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n371_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n402_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT97), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT19), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n336_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n436_));
  AOI211_X1 g235(.A(KEYINPUT108), .B(new_n434_), .C1(new_n402_), .C2(new_n430_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n422_), .A2(new_n424_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n337_), .B1(new_n439_), .B2(new_n373_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n385_), .A2(new_n396_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT99), .B1(new_n373_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT99), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n429_), .A2(new_n444_), .A3(new_n441_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n434_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n335_), .B1(new_n438_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n362_), .A2(new_n372_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n448_), .A2(new_n422_), .A3(new_n424_), .A4(new_n426_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n443_), .A2(new_n445_), .A3(KEYINPUT20), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n435_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n426_), .B(new_n442_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT100), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n435_), .A2(new_n337_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT100), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n448_), .A2(new_n455_), .A3(new_n426_), .A4(new_n442_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n430_), .A2(new_n453_), .A3(new_n454_), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n335_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT27), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT109), .B1(new_n447_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT27), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n430_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n454_), .A2(new_n463_), .B1(new_n450_), .B2(new_n435_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n464_), .B2(new_n335_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n400_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n398_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT20), .B1(new_n429_), .B2(new_n467_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n448_), .A2(new_n426_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n435_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT108), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n431_), .A2(new_n336_), .A3(new_n435_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n446_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n459_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT109), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n465_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n461_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n464_), .A2(new_n335_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n458_), .A2(new_n459_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n462_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT102), .ZN(new_n483_));
  INV_X1    g282(.A(G127gat), .ZN(new_n484_));
  INV_X1    g283(.A(G134gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G113gat), .ZN(new_n487_));
  INV_X1    g286(.A(G120gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G127gat), .A2(G134gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G113gat), .A2(G120gat), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(new_n489_), .A3(new_n490_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n486_), .A2(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n492_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n494_), .B1(KEYINPUT85), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G141gat), .A2(G148gat), .ZN(new_n500_));
  INV_X1    g299(.A(G141gat), .ZN(new_n501_));
  INV_X1    g300(.A(G148gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G155gat), .A2(G162gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(KEYINPUT1), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT1), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n507_), .A2(KEYINPUT87), .A3(G155gat), .A4(G162gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G155gat), .ZN(new_n510_));
  INV_X1    g309(.A(G162gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT86), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(KEYINPUT1), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT86), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(G155gat), .B2(G162gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n500_), .B(new_n503_), .C1(new_n509_), .C2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT3), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n518_), .A2(new_n501_), .A3(new_n502_), .A4(KEYINPUT88), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n520_));
  OAI22_X1  g319(.A1(new_n520_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT2), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n500_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n525_), .A2(new_n512_), .A3(new_n515_), .A4(new_n505_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n499_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n517_), .A2(new_n526_), .A3(new_n498_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n483_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(new_n483_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT4), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G225gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT103), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT4), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n530_), .A2(new_n531_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT104), .B(KEYINPUT0), .Z(new_n542_));
  XNOR2_X1  g341(.A(G1gat), .B(G29gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G85gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n541_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G78gat), .B(G106gat), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n527_), .A2(KEYINPUT29), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n429_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n429_), .A2(KEYINPUT90), .ZN(new_n553_));
  INV_X1    g352(.A(G233gat), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT91), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT91), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(G228gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n557_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n429_), .B(new_n551_), .C1(KEYINPUT90), .C2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n550_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(new_n560_), .A3(new_n550_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n527_), .A2(KEYINPUT29), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G22gat), .B(G50gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n565_), .B(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n561_), .B2(KEYINPUT96), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n562_), .A2(KEYINPUT96), .A3(new_n563_), .A4(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G227gat), .A2(G233gat), .ZN(new_n575_));
  INV_X1    g374(.A(G15gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n499_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT84), .B(G43gat), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G71gat), .B(G99gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n582_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n439_), .A2(KEYINPUT31), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n425_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT30), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n585_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n574_), .A2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n482_), .A2(new_n548_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n548_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n465_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n475_), .B1(new_n465_), .B2(new_n474_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n481_), .B(new_n595_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT110), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n541_), .A2(KEYINPUT33), .A3(new_n547_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT105), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT33), .B1(new_n541_), .B2(new_n547_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n538_), .A2(new_n539_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n532_), .A2(new_n536_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n546_), .B1(new_n607_), .B2(new_n534_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n601_), .A2(new_n602_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n604_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n548_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n451_), .A2(KEYINPUT106), .A3(new_n457_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n438_), .A2(new_n612_), .A3(new_n614_), .A4(new_n446_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n613_), .B1(new_n458_), .B2(KEYINPUT106), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n611_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n574_), .B1(new_n610_), .B2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n477_), .A2(KEYINPUT110), .A3(new_n481_), .A4(new_n595_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n600_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n592_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n594_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT34), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n297_), .A2(new_n237_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n315_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n313_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n237_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n625_), .B(new_n626_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n316_), .A2(new_n237_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n633_), .A2(KEYINPUT35), .A3(new_n624_), .A4(new_n626_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(G134gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(new_n511_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n638_), .B(KEYINPUT36), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n643_), .A3(new_n634_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n307_), .B(new_n649_), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(new_n244_), .ZN(new_n651_));
  XOR2_X1   g450(.A(G183gat), .B(G211gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(G127gat), .B(G155gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT67), .B1(new_n656_), .B2(KEYINPUT17), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n651_), .B(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n656_), .A2(KEYINPUT17), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n641_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n648_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n330_), .A2(new_n622_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n298_), .A3(new_n548_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT38), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n330_), .A2(new_n622_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n660_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n645_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n611_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(G1324gat));
  NAND3_X1  g471(.A1(new_n664_), .A2(new_n299_), .A3(new_n482_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n482_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G8gat), .B1(new_n670_), .B2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT39), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT39), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g478(.A1(new_n664_), .A2(new_n576_), .A3(new_n592_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n667_), .A2(new_n592_), .A3(new_n669_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G15gat), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n682_), .A2(KEYINPUT111), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(KEYINPUT111), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(KEYINPUT41), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(new_n683_), .B2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n680_), .B1(new_n685_), .B2(new_n686_), .ZN(G1326gat));
  OAI21_X1  g486(.A(G22gat), .B1(new_n670_), .B2(new_n574_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT42), .ZN(new_n689_));
  INV_X1    g488(.A(G22gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n664_), .A2(new_n690_), .A3(new_n573_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1327gat));
  INV_X1    g491(.A(new_n286_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n329_), .B(new_n668_), .C1(new_n693_), .C2(new_n284_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n620_), .A2(new_n621_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n594_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n648_), .A2(new_n661_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n700_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n622_), .A2(KEYINPUT43), .A3(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n695_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n699_), .A2(new_n696_), .A3(new_n700_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n622_), .B2(new_n702_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(KEYINPUT44), .A3(new_n695_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n706_), .A2(new_n710_), .A3(new_n548_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(KEYINPUT112), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(KEYINPUT112), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(G29gat), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n645_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n660_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n667_), .A2(new_n716_), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n717_), .A2(G29gat), .A3(new_n611_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT113), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n714_), .A2(new_n721_), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n667_), .A2(new_n724_), .A3(new_n716_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n674_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(new_n674_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT44), .B1(new_n709_), .B2(new_n695_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n705_), .B(new_n694_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n674_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT114), .B1(new_n732_), .B2(new_n724_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n706_), .A2(new_n710_), .A3(new_n482_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(G36gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n729_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n737_), .A2(KEYINPUT115), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n729_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n734_), .A2(new_n735_), .A3(G36gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n735_), .B1(new_n734_), .B2(G36gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT46), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n739_), .A2(new_n745_), .ZN(G1329gat));
  NOR3_X1   g545(.A1(new_n717_), .A2(G43gat), .A3(new_n621_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n706_), .A2(new_n710_), .A3(new_n592_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G43gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g549(.A1(new_n730_), .A2(new_n731_), .A3(new_n574_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n573_), .A2(new_n295_), .ZN(new_n752_));
  OAI22_X1  g551(.A1(new_n751_), .A2(new_n295_), .B1(new_n717_), .B2(new_n752_), .ZN(G1331gat));
  NOR2_X1   g552(.A1(new_n693_), .A2(new_n284_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n329_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n756_), .A2(new_n622_), .A3(new_n663_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n548_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n622_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n669_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n548_), .A2(G57gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n758_), .B1(new_n763_), .B2(new_n764_), .ZN(G1332gat));
  INV_X1    g564(.A(G64gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n757_), .A2(new_n766_), .A3(new_n482_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G64gat), .B1(new_n762_), .B2(new_n674_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n757_), .A2(new_n772_), .A3(new_n592_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G71gat), .B1(new_n762_), .B2(new_n621_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n773_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  NOR2_X1   g576(.A1(new_n574_), .A2(G78gat), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT117), .Z(new_n779_));
  NAND2_X1  g578(.A1(new_n757_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G78gat), .B1(new_n762_), .B2(new_n574_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT50), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT50), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n782_), .B2(new_n783_), .ZN(G1335gat));
  AND2_X1   g583(.A1(new_n759_), .A2(new_n716_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n548_), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n660_), .B(new_n756_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n611_), .A2(new_n213_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(G1336gat));
  AOI21_X1  g588(.A(G92gat), .B1(new_n785_), .B2(new_n482_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n674_), .A2(new_n214_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n787_), .B2(new_n791_), .ZN(G1337gat));
  NAND2_X1  g591(.A1(new_n787_), .A2(new_n592_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n592_), .A2(new_n216_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n793_), .A2(G99gat), .B1(new_n785_), .B2(new_n794_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g595(.A1(new_n785_), .A2(new_n217_), .A3(new_n573_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n787_), .A2(new_n573_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G106gat), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT52), .B(new_n217_), .C1(new_n787_), .C2(new_n573_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n329_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n662_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n805_), .B2(new_n662_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n804_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n809_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT54), .A3(new_n807_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n309_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n325_), .B(new_n816_), .C1(new_n311_), .C2(new_n319_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n328_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n279_), .B2(new_n277_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n267_), .B2(new_n251_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT119), .ZN(new_n822_));
  OR3_X1    g621(.A1(new_n267_), .A2(new_n820_), .A3(new_n251_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n267_), .A2(new_n251_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n820_), .C1(new_n267_), .C2(new_n251_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .A4(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(KEYINPUT120), .A3(new_n828_), .A4(new_n259_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(new_n329_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n827_), .A2(new_n259_), .B1(KEYINPUT120), .B2(new_n828_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n277_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n819_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n815_), .B1(new_n834_), .B2(new_n645_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT58), .ZN(new_n837_));
  INV_X1    g636(.A(new_n818_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n827_), .A2(new_n259_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n828_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n827_), .A2(new_n259_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n277_), .B1(new_n841_), .B2(KEYINPUT56), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n837_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n832_), .B1(new_n839_), .B2(new_n828_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n837_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n818_), .B1(new_n841_), .B2(KEYINPUT56), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n700_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n835_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n829_), .A2(new_n329_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n852_), .A2(new_n832_), .A3(new_n831_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT57), .B(new_n715_), .C1(new_n853_), .C2(new_n819_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n835_), .A2(new_n848_), .A3(KEYINPUT122), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n814_), .B1(new_n856_), .B2(new_n668_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n482_), .A2(new_n593_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n548_), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n857_), .A2(KEYINPUT123), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n835_), .A2(new_n854_), .A3(new_n848_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n862_), .A2(new_n668_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n611_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n858_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT59), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT123), .B1(new_n857_), .B2(new_n860_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n755_), .A2(new_n487_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n861_), .A2(new_n866_), .A3(new_n867_), .A4(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n487_), .B1(new_n865_), .B2(new_n755_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1340gat));
  INV_X1    g670(.A(new_n865_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n488_), .B1(new_n287_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n872_), .B(new_n873_), .C1(KEYINPUT60), .C2(new_n488_), .ZN(new_n874_));
  AND4_X1   g673(.A1(new_n754_), .A2(new_n861_), .A3(new_n866_), .A4(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n488_), .ZN(G1341gat));
  NOR2_X1   g675(.A1(new_n668_), .A2(new_n484_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n861_), .A2(new_n866_), .A3(new_n867_), .A4(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n484_), .B1(new_n865_), .B2(new_n668_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1342gat));
  NOR2_X1   g679(.A1(new_n702_), .A2(new_n485_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n861_), .A2(new_n866_), .A3(new_n867_), .A4(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n485_), .B1(new_n865_), .B2(new_n715_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1343gat));
  NOR3_X1   g683(.A1(new_n863_), .A2(new_n611_), .A3(new_n592_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n674_), .A2(new_n573_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n755_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n501_), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n287_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n502_), .ZN(G1345gat));
  NOR2_X1   g691(.A1(new_n888_), .A2(new_n668_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT61), .B(G155gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  OAI21_X1  g694(.A(new_n511_), .B1(new_n888_), .B2(new_n715_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n700_), .A2(G162gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT124), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n885_), .A2(new_n887_), .A3(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n674_), .A2(new_n548_), .A3(new_n593_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n857_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n329_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G169gat), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n907_), .B(new_n908_), .C1(new_n384_), .C2(new_n904_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n903_), .B2(new_n754_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n863_), .A2(new_n902_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n287_), .A2(new_n413_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  AOI21_X1  g712(.A(G183gat), .B1(new_n911_), .B2(new_n660_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n668_), .A2(new_n391_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n903_), .B2(new_n915_), .ZN(G1350gat));
  INV_X1    g715(.A(new_n903_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G190gat), .B1(new_n917_), .B2(new_n702_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n903_), .A2(new_n390_), .A3(new_n645_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1351gat));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n862_), .A2(new_n668_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n592_), .B1(new_n922_), .B2(new_n813_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n482_), .A2(new_n595_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n921_), .B1(new_n923_), .B2(new_n925_), .ZN(new_n926_));
  NOR4_X1   g725(.A1(new_n863_), .A2(KEYINPUT125), .A3(new_n592_), .A4(new_n924_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n329_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g729(.A1(new_n258_), .A2(KEYINPUT126), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n928_), .B2(new_n754_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n928_), .A2(new_n754_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n368_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1353gat));
  OR2_X1    g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n936_), .B1(new_n928_), .B2(new_n660_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n928_), .A2(new_n660_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT63), .B(G211gat), .Z(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(G1354gat));
  OAI21_X1  g739(.A(new_n645_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT127), .ZN(new_n942_));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n944_), .B(new_n645_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n943_), .A3(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n928_), .A2(G218gat), .A3(new_n700_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1355gat));
endmodule


