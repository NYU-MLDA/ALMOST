//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT72), .B(G8gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G1gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT73), .B1(new_n205_), .B2(KEYINPUT14), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208_));
  AOI211_X1 g007(.A(new_n207_), .B(new_n208_), .C1(new_n204_), .C2(G1gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n203_), .B1(new_n206_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n203_), .B(new_n211_), .C1(new_n206_), .C2(new_n209_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G29gat), .B(G36gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n219_), .B(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(KEYINPUT78), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT78), .B1(new_n215_), .B2(new_n223_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n202_), .B(new_n221_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n215_), .A2(new_n223_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n223_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n231_), .A2(new_n213_), .A3(KEYINPUT79), .A4(new_n214_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n215_), .B2(new_n223_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n230_), .A2(new_n224_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n227_), .B1(new_n235_), .B2(new_n202_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G113gat), .B(G141gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT80), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n227_), .B(new_n240_), .C1(new_n235_), .C2(new_n202_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT23), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(KEYINPUT83), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(KEYINPUT23), .ZN(new_n249_));
  NOR3_X1   g048(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(G169gat), .B2(G176gat), .ZN(new_n252_));
  INV_X1    g051(.A(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(G176gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT82), .B(G190gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(KEYINPUT26), .ZN(new_n259_));
  INV_X1    g058(.A(G183gat), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(KEYINPUT25), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT81), .ZN(new_n262_));
  OR3_X1    g061(.A1(new_n260_), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(KEYINPUT25), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n249_), .B(new_n256_), .C1(new_n259_), .C2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G169gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n246_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n248_), .B2(new_n269_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n258_), .A2(G183gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(G15gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT30), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n274_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G113gat), .B(G120gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n279_), .B(new_n280_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n284_), .B2(new_n282_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n278_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287_));
  INV_X1    g086(.A(G43gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT31), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n290_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT26), .B(G190gat), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n261_), .A2(new_n264_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n256_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(new_n271_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n253_), .A2(new_n254_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT22), .B(G169gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT90), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n302_), .B2(new_n254_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n249_), .B1(G183gat), .B2(G190gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n299_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307_));
  INV_X1    g106(.A(G204gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G197gat), .ZN(new_n309_));
  INV_X1    g108(.A(G197gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G204gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT87), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT21), .B1(new_n309_), .B2(KEYINPUT87), .ZN(new_n315_));
  OAI221_X1 g114(.A(new_n307_), .B1(new_n312_), .B2(new_n313_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(KEYINPUT21), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n317_), .A2(new_n307_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n295_), .B1(new_n306_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n316_), .A2(new_n318_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n273_), .A3(new_n266_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n303_), .A2(new_n304_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n299_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n325_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n274_), .A2(new_n319_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT20), .ZN(new_n332_));
  INV_X1    g131(.A(new_n324_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT94), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n326_), .B(KEYINPUT20), .C1(new_n325_), .C2(new_n305_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n327_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n335_), .B2(new_n333_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT20), .A4(new_n324_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n335_), .A2(new_n345_), .A3(new_n333_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .A4(new_n342_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(KEYINPUT1), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n353_), .B2(KEYINPUT1), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n354_), .B2(KEYINPUT85), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT85), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n356_), .B(new_n351_), .C1(new_n353_), .C2(KEYINPUT1), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G141gat), .B(G148gat), .Z(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT86), .ZN(new_n362_));
  NOR3_X1   g161(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n363_));
  AND3_X1   g162(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n351_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(new_n353_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n360_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n285_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n360_), .A2(new_n370_), .A3(new_n284_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT92), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n371_), .A2(new_n378_), .A3(new_n285_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT93), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT4), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n381_), .A2(new_n376_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n377_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  AOI211_X1 g188(.A(new_n377_), .B(new_n387_), .C1(new_n380_), .C2(new_n382_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n344_), .B(new_n350_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n381_), .A2(new_n376_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n379_), .A2(KEYINPUT93), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n379_), .A2(KEYINPUT93), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NOR4_X1   g194(.A1(new_n395_), .A2(KEYINPUT33), .A3(new_n377_), .A4(new_n387_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n347_), .A2(new_n341_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n341_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n349_), .A2(new_n348_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(new_n346_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n376_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n380_), .A2(new_n404_), .A3(new_n381_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n405_), .B(new_n387_), .C1(new_n374_), .C2(new_n404_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n400_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n391_), .B1(new_n399_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT28), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n319_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n410_), .A2(new_n412_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(G78gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G106gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G22gat), .B(G50gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OR3_X1    g221(.A1(new_n413_), .A2(new_n414_), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n408_), .A2(KEYINPUT95), .A3(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n389_), .A2(new_n390_), .A3(KEYINPUT96), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n387_), .B1(new_n395_), .B2(new_n377_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n383_), .A2(new_n388_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n337_), .A2(new_n401_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT97), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT97), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n337_), .A2(new_n436_), .A3(new_n401_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n435_), .A2(KEYINPUT27), .A3(new_n400_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n403_), .A2(new_n400_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT27), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n433_), .A2(new_n438_), .A3(new_n441_), .A4(new_n425_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n427_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT95), .B1(new_n408_), .B2(new_n426_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n294_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n433_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(new_n294_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n438_), .A2(new_n441_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n448_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n447_), .B(new_n426_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n245_), .B1(new_n445_), .B2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G85gat), .A2(G92gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n418_), .A4(KEYINPUT66), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n462_));
  OAI22_X1  g261(.A1(new_n462_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT67), .B(new_n455_), .C1(new_n458_), .C2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT68), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n453_), .A2(new_n454_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n458_), .B1(new_n469_), .B2(KEYINPUT9), .ZN(new_n470_));
  OR2_X1    g269(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT64), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n418_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n454_), .A2(KEYINPUT9), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n470_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n465_), .A2(KEYINPUT68), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(new_n455_), .C1(new_n458_), .C2(new_n464_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT8), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n467_), .B(new_n479_), .C1(new_n480_), .C2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G57gat), .B(G64gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n486_));
  XOR2_X1   g285(.A(G71gat), .B(G78gat), .Z(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT12), .B1(new_n484_), .B2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n484_), .A2(new_n492_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT69), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n483_), .B1(KEYINPUT68), .B2(new_n465_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n467_), .A2(new_n479_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n465_), .A2(KEYINPUT68), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT8), .A3(new_n482_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n502_), .A2(KEYINPUT69), .A3(new_n467_), .A4(new_n479_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n492_), .A2(KEYINPUT12), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n495_), .A2(new_n496_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n496_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n499_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n491_), .B1(new_n509_), .B2(new_n502_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n510_), .B2(new_n494_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G120gat), .B(G148gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT5), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G176gat), .B(G204gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n512_), .B(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT13), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT13), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(G231gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n491_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n216_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G127gat), .B(G155gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G183gat), .B(G211gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n524_), .A2(KEYINPUT75), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT75), .B1(new_n524_), .B2(new_n531_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n529_), .B(new_n530_), .ZN(new_n534_));
  OAI22_X1  g333(.A1(new_n532_), .A2(new_n533_), .B1(new_n524_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT76), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n500_), .A2(new_n220_), .A3(new_n503_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT35), .ZN(new_n542_));
  INV_X1    g341(.A(new_n484_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(new_n219_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(KEYINPUT35), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT71), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n538_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n544_), .B2(new_n538_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n553_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n521_), .A2(new_n537_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n452_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT99), .ZN(new_n564_));
  INV_X1    g363(.A(G1gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n446_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT38), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n556_), .A2(new_n558_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT100), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n556_), .A2(new_n571_), .A3(new_n558_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n445_), .B2(new_n451_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n521_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n244_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(new_n535_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n580_), .B2(new_n433_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n566_), .A2(new_n567_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n568_), .A2(new_n581_), .A3(new_n582_), .ZN(G1324gat));
  NOR2_X1   g382(.A1(new_n449_), .A2(new_n450_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n204_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n564_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n579_), .A2(new_n584_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n589_));
  AND4_X1   g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .A4(G8gat), .ZN(new_n590_));
  INV_X1    g389(.A(G8gat), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(KEYINPUT101), .B2(KEYINPUT39), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n588_), .A2(new_n592_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n586_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g394(.A(KEYINPUT41), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n579_), .A2(new_n293_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(G15gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n597_), .B2(G15gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n596_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(KEYINPUT41), .A3(new_n599_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n563_), .A2(G15gat), .A3(new_n294_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT103), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n602_), .A2(new_n604_), .A3(new_n608_), .A4(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(G1326gat));
  OAI21_X1  g409(.A(G22gat), .B1(new_n580_), .B2(new_n426_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT42), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n426_), .A2(G22gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n563_), .B2(new_n613_), .ZN(G1327gat));
  NOR2_X1   g413(.A1(new_n577_), .A2(new_n536_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n445_), .A2(new_n451_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n617_), .B2(new_n561_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n561_), .ZN(new_n619_));
  AOI211_X1 g418(.A(KEYINPUT43), .B(new_n619_), .C1(new_n445_), .C2(new_n451_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n615_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT44), .B(new_n615_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n446_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(G29gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n574_), .A2(KEYINPUT104), .A3(new_n537_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n536_), .B2(new_n573_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n521_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n452_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n433_), .A2(G29gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT105), .Z(new_n634_));
  OAI21_X1  g433(.A(new_n627_), .B1(new_n632_), .B2(new_n634_), .ZN(G1328gat));
  NOR2_X1   g434(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT107), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n623_), .A2(new_n584_), .A3(new_n624_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G36gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n584_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n632_), .A2(G36gat), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT45), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n637_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n645_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n637_), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n647_), .B(new_n648_), .C1(new_n639_), .C2(new_n643_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1329gat));
  NAND3_X1  g449(.A1(new_n625_), .A2(G43gat), .A3(new_n293_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n288_), .B1(new_n632_), .B2(new_n294_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT108), .Z(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT47), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT47), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n651_), .A2(new_n656_), .A3(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1330gat));
  OR3_X1    g457(.A1(new_n632_), .A2(G50gat), .A3(new_n426_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n625_), .A2(new_n660_), .A3(new_n425_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G50gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n625_), .B2(new_n425_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1331gat));
  AOI21_X1  g463(.A(new_n244_), .B1(new_n445_), .B2(new_n451_), .ZN(new_n665_));
  AND4_X1   g464(.A1(new_n521_), .A2(new_n665_), .A3(new_n536_), .A4(new_n619_), .ZN(new_n666_));
  INV_X1    g465(.A(G57gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n446_), .ZN(new_n668_));
  AND4_X1   g467(.A1(new_n245_), .A2(new_n575_), .A3(new_n521_), .A4(new_n536_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(new_n446_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n670_), .B2(new_n667_), .ZN(G1332gat));
  INV_X1    g470(.A(G64gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n669_), .B2(new_n584_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT48), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n584_), .A2(new_n672_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT110), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n666_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(G1333gat));
  INV_X1    g477(.A(G71gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n669_), .B2(new_n293_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT49), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n666_), .A2(new_n679_), .A3(new_n293_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1334gat));
  AOI21_X1  g482(.A(new_n416_), .B1(new_n669_), .B2(new_n425_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT50), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n666_), .A2(new_n416_), .A3(new_n425_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1335gat));
  OR2_X1    g486(.A1(new_n618_), .A2(new_n620_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n576_), .A2(new_n244_), .A3(new_n536_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G85gat), .B1(new_n690_), .B2(new_n433_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n576_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n665_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G85gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n446_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1336gat));
  AOI21_X1  g495(.A(G92gat), .B1(new_n693_), .B2(new_n584_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n690_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n584_), .A2(G92gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT111), .Z(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n698_), .B2(new_n700_), .ZN(G1337gat));
  OAI21_X1  g500(.A(G99gat), .B1(new_n690_), .B2(new_n294_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT112), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n693_), .B(new_n293_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g505(.A1(new_n693_), .A2(new_n418_), .A3(new_n425_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n425_), .B(new_n689_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT52), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G106gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G106gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g512(.A1(new_n507_), .A2(new_n511_), .A3(new_n517_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n244_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n509_), .A2(new_n491_), .A3(new_n502_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n484_), .A2(new_n492_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT12), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AND4_X1   g518(.A1(new_n496_), .A2(new_n506_), .A3(new_n716_), .A4(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n506_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n510_), .B2(KEYINPUT12), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n508_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(KEYINPUT55), .B2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n495_), .A2(KEYINPUT55), .A3(new_n496_), .A4(new_n506_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n516_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT113), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n496_), .B1(new_n495_), .B2(new_n506_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n507_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n517_), .B1(new_n734_), .B2(new_n725_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n729_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n715_), .B1(new_n731_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n202_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(new_n221_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n739_), .B(new_n241_), .C1(new_n235_), .C2(new_n738_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n243_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n518_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n573_), .B1(new_n737_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT57), .B(new_n573_), .C1(new_n737_), .C2(new_n742_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT58), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n243_), .A2(new_n740_), .A3(new_n714_), .ZN(new_n748_));
  AND2_X1   g547(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n735_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n749_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n517_), .B(new_n754_), .C1(new_n734_), .C2(new_n725_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n747_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(KEYINPUT115), .A3(new_n561_), .ZN(new_n757_));
  OR3_X1    g556(.A1(new_n751_), .A2(new_n747_), .A3(new_n755_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT115), .B1(new_n756_), .B2(new_n561_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n745_), .B(new_n746_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n756_), .A2(new_n561_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n758_), .A3(new_n757_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(KEYINPUT116), .A3(new_n745_), .A4(new_n746_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n763_), .A2(new_n535_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n562_), .A2(new_n245_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT54), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NOR4_X1   g571(.A1(new_n584_), .A2(new_n425_), .A3(new_n433_), .A4(new_n294_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n244_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(KEYINPUT59), .ZN(new_n777_));
  INV_X1    g576(.A(new_n761_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n771_), .B1(new_n536_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n773_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n244_), .A2(G113gat), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT117), .Z(new_n785_));
  AOI21_X1  g584(.A(new_n776_), .B1(new_n783_), .B2(new_n785_), .ZN(G1340gat));
  OAI21_X1  g585(.A(G120gat), .B1(new_n782_), .B2(new_n576_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n788_));
  AOI21_X1  g587(.A(G120gat), .B1(new_n521_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n788_), .B2(G120gat), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n775_), .A2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT118), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(KEYINPUT118), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n787_), .B1(new_n792_), .B2(new_n793_), .ZN(G1341gat));
  INV_X1    g593(.A(G127gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n774_), .B2(new_n537_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n797_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n535_), .A2(new_n795_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n798_), .A2(new_n799_), .B1(new_n783_), .B2(new_n800_), .ZN(G1342gat));
  INV_X1    g600(.A(G134gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n619_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n774_), .B2(new_n573_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT120), .B(new_n802_), .C1(new_n774_), .C2(new_n573_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n783_), .A2(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(G1343gat));
  NOR4_X1   g607(.A1(new_n584_), .A2(new_n426_), .A3(new_n433_), .A4(new_n293_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n772_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n244_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n521_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g614(.A1(new_n810_), .A2(new_n537_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT61), .B(G155gat), .Z(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1346gat));
  AOI21_X1  g617(.A(G162gat), .B1(new_n811_), .B2(new_n574_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n561_), .A2(G162gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT121), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n811_), .B2(new_n821_), .ZN(G1347gat));
  NAND2_X1  g621(.A1(new_n584_), .A2(new_n447_), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT122), .Z(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n425_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n779_), .A2(new_n244_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT62), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n826_), .A2(new_n827_), .A3(G169gat), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n779_), .A2(new_n302_), .A3(new_n244_), .A4(new_n825_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n826_), .B2(G169gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(G1348gat));
  NAND2_X1  g630(.A1(new_n779_), .A2(new_n825_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n254_), .B1(new_n832_), .B2(new_n576_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT123), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(KEYINPUT123), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n772_), .A2(new_n426_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n824_), .A2(new_n254_), .A3(new_n576_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n834_), .A2(new_n835_), .B1(new_n837_), .B2(new_n838_), .ZN(G1349gat));
  AOI211_X1 g638(.A(new_n535_), .B(new_n832_), .C1(new_n261_), .C2(new_n264_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n836_), .A2(new_n537_), .A3(new_n824_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n841_), .A2(KEYINPUT124), .ZN(new_n842_));
  AOI21_X1  g641(.A(G183gat), .B1(new_n841_), .B2(KEYINPUT124), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n840_), .B1(new_n842_), .B2(new_n843_), .ZN(G1350gat));
  OR3_X1    g643(.A1(new_n832_), .A2(new_n296_), .A3(new_n573_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G190gat), .B1(new_n832_), .B2(new_n619_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(KEYINPUT125), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(KEYINPUT125), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n847_), .B2(new_n848_), .ZN(G1351gat));
  NOR2_X1   g648(.A1(new_n446_), .A2(new_n426_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n584_), .A2(new_n294_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n244_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n521_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g655(.A(new_n535_), .B(new_n851_), .C1(new_n769_), .C2(new_n771_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT63), .B(G211gat), .Z(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n857_), .B2(new_n859_), .ZN(G1354gat));
  NAND3_X1  g659(.A1(new_n852_), .A2(G218gat), .A3(new_n561_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT126), .ZN(new_n862_));
  INV_X1    g661(.A(new_n851_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n772_), .A2(new_n862_), .A3(new_n574_), .A4(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(G218gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n862_), .B1(new_n852_), .B2(new_n574_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n861_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT127), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT127), .B(new_n861_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1355gat));
endmodule


