//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT16), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G183gat), .B(G211gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT17), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n208_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n211_), .A2(new_n212_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G1gat), .B(G8gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n215_), .B(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G57gat), .B(G64gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n220_));
  XOR2_X1   g019(.A(G71gat), .B(G78gat), .Z(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n220_), .A2(new_n221_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n218_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G231gat), .A2(G233gat), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n228_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n207_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n205_), .A2(new_n206_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G169gat), .B(G197gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT77), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT71), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n241_), .A2(KEYINPUT71), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(KEYINPUT71), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT15), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n218_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G229gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(new_n218_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT76), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n251_), .A2(new_n258_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n253_), .B(new_n218_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n252_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n240_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n263_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n239_), .A3(new_n256_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(G169gat), .B2(G176gat), .ZN(new_n272_));
  INV_X1    g071(.A(G169gat), .ZN(new_n273_));
  INV_X1    g072(.A(G176gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n270_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT23), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G183gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT25), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT78), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G190gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT25), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G183gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT79), .B1(new_n285_), .B2(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT78), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n282_), .A3(KEYINPUT25), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT79), .ZN(new_n293_));
  INV_X1    g092(.A(G190gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT26), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n276_), .B(new_n281_), .C1(new_n289_), .C2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n277_), .A2(new_n299_), .A3(KEYINPUT23), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n277_), .B2(KEYINPUT23), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n280_), .A2(KEYINPUT82), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n304_), .A2(new_n279_), .A3(G183gat), .A4(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n298_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n273_), .A2(new_n274_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n274_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n273_), .A2(KEYINPUT22), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n309_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n297_), .B1(new_n307_), .B2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT30), .Z(new_n319_));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G15gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT83), .B(G43gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n321_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n319_), .A2(new_n320_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n321_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G134gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G127gat), .ZN(new_n333_));
  INV_X1    g132(.A(G127gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G134gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G120gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G113gat), .ZN(new_n338_));
  INV_X1    g137(.A(G113gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G120gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n333_), .A2(new_n335_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(KEYINPUT85), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n336_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT31), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n331_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n328_), .A2(new_n330_), .A3(new_n349_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  INV_X1    g153(.A(G141gat), .ZN(new_n355_));
  INV_X1    g154(.A(G148gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT2), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n355_), .A2(new_n356_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .A4(new_n358_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n380_));
  INV_X1    g179(.A(G204gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(G197gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(G197gat), .ZN(new_n383_));
  INV_X1    g182(.A(G197gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n379_), .A2(new_n386_), .A3(KEYINPUT21), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(G204gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n383_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT21), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n378_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n386_), .A2(KEYINPUT21), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n387_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n377_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G78gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n397_), .A2(G78gat), .ZN(new_n400_));
  INV_X1    g199(.A(G106gat), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n397_), .A2(G78gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(G106gat), .B1(new_n403_), .B2(new_n398_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n376_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n401_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(G106gat), .A3(new_n398_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n376_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n394_), .A2(new_n395_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G22gat), .B(G50gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n411_), .B(new_n412_), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n405_), .A2(new_n413_), .A3(new_n409_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT97), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n344_), .A2(new_n347_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n342_), .A2(new_n343_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n420_), .A2(new_n372_), .A3(new_n367_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n418_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n348_), .A2(new_n373_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT97), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n422_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G85gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT98), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT98), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(new_n436_), .A3(new_n433_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT95), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n423_), .B2(KEYINPUT4), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n419_), .A2(KEYINPUT95), .A3(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n419_), .A2(new_n421_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n439_), .A2(new_n441_), .B1(new_n442_), .B2(KEYINPUT4), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n426_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n435_), .A2(new_n437_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT99), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n434_), .A2(KEYINPUT98), .B1(new_n443_), .B2(new_n426_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT99), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n437_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n423_), .A2(KEYINPUT4), .A3(new_n424_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n441_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT95), .B1(new_n419_), .B2(new_n440_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n427_), .B(new_n450_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n442_), .A2(new_n426_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n432_), .ZN(new_n455_));
  OR2_X1    g254(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n446_), .A2(new_n449_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n461_));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT94), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n462_), .A2(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n461_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n461_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n464_), .A3(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G8gat), .B(G36gat), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n467_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT20), .B1(new_n318_), .B2(new_n393_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n311_), .A2(new_n315_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n309_), .B1(new_n478_), .B2(G176gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT91), .B(new_n309_), .C1(new_n478_), .C2(G176gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n298_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n281_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n283_), .A2(new_n288_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n294_), .A2(KEYINPUT26), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n488_), .A2(new_n286_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n488_), .B2(new_n286_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n487_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n272_), .A2(new_n275_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(KEYINPUT90), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n270_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT90), .B1(new_n492_), .B2(new_n493_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n485_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n477_), .B1(new_n498_), .B2(new_n393_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G226gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT19), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n476_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n393_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n285_), .A2(G190gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n294_), .A2(KEYINPUT26), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT89), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n488_), .A2(new_n286_), .A3(new_n489_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n486_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n493_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n505_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n504_), .B1(new_n513_), .B2(new_n485_), .ZN(new_n514_));
  OAI211_X1 g313(.A(KEYINPUT92), .B(new_n501_), .C1(new_n514_), .C2(new_n477_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n503_), .A2(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n504_), .B(new_n485_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n318_), .B2(new_n393_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n502_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n475_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  AOI211_X1 g321(.A(new_n522_), .B(new_n474_), .C1(new_n503_), .C2(new_n515_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT102), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT32), .B1(new_n472_), .B2(new_n473_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n477_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n485_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n270_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n303_), .A2(new_n305_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n278_), .A2(KEYINPUT81), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n277_), .A2(new_n299_), .A3(KEYINPUT23), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n530_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n508_), .A2(new_n509_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n511_), .B1(new_n536_), .B2(new_n487_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n537_), .B2(KEYINPUT90), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n529_), .B1(new_n538_), .B2(new_n512_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n528_), .B(new_n502_), .C1(new_n539_), .C2(new_n504_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT101), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n502_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n542_), .A2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n527_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n526_), .A2(KEYINPUT100), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT100), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n547_), .B(KEYINPUT32), .C1(new_n472_), .C2(new_n473_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n546_), .A2(new_n520_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n528_), .B1(new_n539_), .B2(new_n504_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT92), .B1(new_n550_), .B2(new_n501_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n515_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n453_), .A2(new_n454_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n433_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n455_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n545_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n460_), .A2(new_n524_), .B1(new_n525_), .B2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n545_), .A2(new_n553_), .A3(new_n556_), .A4(KEYINPUT102), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n417_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT27), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n556_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n516_), .A2(new_n520_), .A3(new_n475_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n474_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(KEYINPUT27), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n562_), .A2(new_n417_), .A3(new_n563_), .A4(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n353_), .B1(new_n560_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT103), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n520_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n474_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT27), .B1(new_n572_), .B2(new_n564_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n564_), .A2(KEYINPUT27), .A3(new_n565_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n570_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n562_), .A2(KEYINPUT103), .A3(new_n566_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n417_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n353_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n577_), .A2(new_n563_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n269_), .B1(new_n569_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT6), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT10), .B(G99gat), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n401_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G85gat), .B(G92gat), .Z(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT9), .ZN(new_n590_));
  INV_X1    g389(.A(G85gat), .ZN(new_n591_));
  INV_X1    g390(.A(G92gat), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT9), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n586_), .A2(new_n588_), .A3(new_n590_), .A4(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT7), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n589_), .B1(new_n597_), .B2(new_n585_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n598_), .A2(KEYINPUT8), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(KEYINPUT8), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n594_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT65), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(KEYINPUT12), .A3(new_n225_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT64), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n225_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n601_), .A2(new_n225_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n608_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n606_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT66), .B(KEYINPUT5), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT67), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n613_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n582_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(KEYINPUT13), .A3(new_n622_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT68), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT74), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n603_), .A2(new_n250_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n633_));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  OAI22_X1  g434(.A1(new_n601_), .A2(new_n253_), .B1(KEYINPUT35), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT35), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT70), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n632_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT73), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n632_), .A2(KEYINPUT73), .A3(new_n639_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT72), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n636_), .A2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n636_), .A2(new_n644_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n632_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n642_), .A2(new_n643_), .B1(new_n638_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G190gat), .B(G218gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT36), .Z(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n631_), .B1(new_n648_), .B2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n651_), .A2(KEYINPUT36), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n632_), .A2(KEYINPUT73), .A3(new_n639_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT73), .B1(new_n632_), .B2(new_n639_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n647_), .A2(new_n638_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT74), .B(new_n652_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n654_), .A2(new_n656_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT37), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n652_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n648_), .B2(new_n655_), .ZN(new_n665_));
  AOI22_X1  g464(.A1(new_n662_), .A2(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  AND4_X1   g465(.A1(new_n234_), .A2(new_n581_), .A3(new_n630_), .A4(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n556_), .B(KEYINPUT104), .Z(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n209_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n662_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n569_), .B2(new_n580_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n234_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n628_), .A2(new_n673_), .A3(new_n269_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n556_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G1gat), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n670_), .ZN(new_n678_));
  MUX2_X1   g477(.A(new_n670_), .B(new_n678_), .S(KEYINPUT38), .Z(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT105), .ZN(G1324gat));
  INV_X1    g479(.A(new_n577_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n675_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G8gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT39), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n667_), .A2(new_n210_), .A3(new_n681_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n684_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n684_), .B2(new_n687_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1325gat));
  INV_X1    g490(.A(G15gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n675_), .B2(new_n579_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT41), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n667_), .A2(new_n692_), .A3(new_n579_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1326gat));
  INV_X1    g495(.A(G22gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n675_), .B2(new_n417_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT42), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n667_), .A2(new_n697_), .A3(new_n417_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n671_), .A2(new_n673_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n628_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n581_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n556_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n666_), .B1(new_n569_), .B2(new_n580_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n706_), .B(KEYINPUT43), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n628_), .A2(new_n234_), .A3(new_n269_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n707_), .B2(new_n706_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n662_), .A2(new_n663_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n665_), .A2(new_n664_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n557_), .A2(new_n525_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n457_), .A2(new_n459_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n449_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n448_), .B1(new_n447_), .B2(new_n437_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n572_), .A2(new_n564_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n716_), .B(new_n559_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n578_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n579_), .B1(new_n723_), .B2(new_n567_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n351_), .A2(new_n415_), .A3(new_n416_), .A4(new_n352_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n556_), .B(new_n725_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n715_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT109), .B1(new_n727_), .B2(KEYINPUT108), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n709_), .B(new_n710_), .C1(new_n712_), .C2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT43), .B1(new_n727_), .B2(KEYINPUT109), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n734_), .A2(KEYINPUT44), .A3(new_n709_), .A4(new_n710_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n669_), .A2(G29gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n705_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  NAND3_X1  g538(.A1(new_n731_), .A2(new_n681_), .A3(new_n735_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G36gat), .ZN(new_n741_));
  INV_X1    g540(.A(G36gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n704_), .A2(new_n742_), .A3(new_n681_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT45), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n741_), .A2(KEYINPUT46), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1329gat));
  XOR2_X1   g548(.A(KEYINPUT110), .B(G43gat), .Z(new_n750_));
  INV_X1    g549(.A(new_n704_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n353_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n579_), .A2(G43gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n736_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g554(.A(G50gat), .B1(new_n704_), .B2(new_n417_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n417_), .A2(G50gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n737_), .B2(new_n757_), .ZN(G1331gat));
  INV_X1    g557(.A(new_n269_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n569_), .B2(new_n580_), .ZN(new_n760_));
  AND4_X1   g559(.A1(new_n234_), .A2(new_n760_), .A3(new_n628_), .A4(new_n666_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n669_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT111), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n234_), .A2(new_n264_), .A3(new_n267_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n629_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n672_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n556_), .A2(G57gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(G1332gat));
  OAI21_X1  g568(.A(G64gat), .B1(new_n766_), .B2(new_n577_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT48), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n577_), .A2(G64gat), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT112), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n761_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(new_n774_), .ZN(G1333gat));
  INV_X1    g574(.A(G71gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n761_), .A2(new_n776_), .A3(new_n579_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n767_), .A2(new_n579_), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(G71gat), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G71gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT114), .ZN(G1334gat));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n761_), .A2(new_n784_), .A3(new_n417_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n767_), .B2(new_n417_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n787_));
  AND2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n786_), .A2(new_n787_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1335gat));
  AND4_X1   g589(.A1(new_n671_), .A2(new_n760_), .A3(new_n673_), .A4(new_n629_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n591_), .A3(new_n669_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n628_), .A2(new_n673_), .A3(new_n269_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n709_), .B1(new_n712_), .B2(new_n728_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT116), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n734_), .A2(new_n796_), .A3(new_n709_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(new_n556_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n792_), .B1(new_n799_), .B2(new_n591_), .ZN(G1336gat));
  AOI21_X1  g599(.A(G92gat), .B1(new_n791_), .B2(new_n681_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT117), .Z(new_n802_));
  NOR2_X1   g601(.A1(new_n577_), .A2(new_n592_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n798_), .B2(new_n803_), .ZN(G1337gat));
  INV_X1    g603(.A(G99gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n798_), .B2(new_n579_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n791_), .A2(new_n587_), .A3(new_n579_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n353_), .B(new_n793_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n810_), .B(new_n807_), .C1(new_n811_), .C2(new_n805_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n791_), .A2(new_n401_), .A3(new_n417_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n401_), .B1(new_n817_), .B2(KEYINPUT52), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n793_), .A2(new_n578_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n794_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(KEYINPUT119), .A3(new_n821_), .ZN(new_n822_));
  OAI221_X1 g621(.A(new_n818_), .B1(new_n817_), .B2(KEYINPUT52), .C1(new_n794_), .C2(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT53), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n816_), .A2(new_n822_), .A3(new_n826_), .A4(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1339gat));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n764_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n830_));
  AND4_X1   g629(.A1(new_n829_), .A2(new_n713_), .A3(new_n714_), .A4(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n666_), .B2(new_n830_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n251_), .A2(new_n254_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n251_), .A2(KEYINPUT121), .A3(new_n254_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n252_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n260_), .A2(new_n261_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n238_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n266_), .A2(new_n237_), .A3(new_n256_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n840_), .B(new_n841_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n613_), .A2(new_n615_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n264_), .A2(new_n267_), .B1(new_n843_), .B2(new_n621_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n607_), .B1(new_n604_), .B2(new_n612_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n613_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n604_), .A2(new_n612_), .A3(KEYINPUT55), .A4(new_n607_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n621_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n844_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n849_), .A2(new_n850_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n842_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n662_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n857_));
  OR3_X1    g656(.A1(new_n849_), .A2(KEYINPUT122), .A3(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n849_), .A2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n840_), .A2(new_n622_), .A3(new_n841_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n858_), .A2(KEYINPUT58), .A3(new_n860_), .A4(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n861_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n849_), .A2(KEYINPUT122), .A3(new_n857_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(new_n715_), .A3(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n853_), .A2(KEYINPUT57), .A3(new_n662_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n856_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n833_), .B1(new_n869_), .B2(new_n673_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n681_), .A2(new_n725_), .A3(new_n668_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n339_), .A3(new_n759_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(KEYINPUT123), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n853_), .A2(KEYINPUT57), .A3(new_n662_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n853_), .B2(new_n662_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n234_), .B1(new_n880_), .B2(new_n867_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n871_), .B(new_n877_), .C1(new_n881_), .C2(new_n833_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n269_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n874_), .B1(new_n888_), .B2(new_n339_), .ZN(G1340gat));
  INV_X1    g688(.A(new_n628_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n337_), .B1(new_n890_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n873_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n337_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n882_), .A2(new_n884_), .A3(new_n629_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n337_), .ZN(G1341gat));
  AOI21_X1  g693(.A(G127gat), .B1(new_n873_), .B2(new_n234_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n886_), .A2(new_n887_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n234_), .A2(G127gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT125), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n896_), .B2(new_n898_), .ZN(G1342gat));
  NAND3_X1  g698(.A1(new_n873_), .A2(new_n332_), .A3(new_n671_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n886_), .A2(new_n887_), .A3(new_n666_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n332_), .ZN(G1343gat));
  NOR2_X1   g701(.A1(new_n870_), .A2(new_n579_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n681_), .A2(new_n578_), .A3(new_n668_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n759_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n629_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n234_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT61), .B(G155gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  AOI21_X1  g711(.A(G162gat), .B1(new_n905_), .B2(new_n671_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n715_), .A2(G162gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT126), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n905_), .B2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  INV_X1    g716(.A(new_n870_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n577_), .A2(new_n725_), .A3(new_n669_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n269_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n917_), .B1(new_n921_), .B2(new_n273_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n923_));
  OAI211_X1 g722(.A(KEYINPUT62), .B(G169gat), .C1(new_n920_), .C2(new_n269_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(G1348gat));
  OAI21_X1  g724(.A(G176gat), .B1(new_n920_), .B2(new_n630_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n628_), .A2(new_n274_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n920_), .B2(new_n927_), .ZN(G1349gat));
  NOR2_X1   g727(.A1(new_n920_), .A2(new_n673_), .ZN(new_n929_));
  MUX2_X1   g728(.A(G183gat), .B(new_n487_), .S(new_n929_), .Z(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n920_), .B2(new_n666_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n671_), .A2(new_n536_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n920_), .B2(new_n932_), .ZN(G1351gat));
  NAND4_X1  g732(.A1(new_n903_), .A2(new_n563_), .A3(new_n417_), .A4(new_n681_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n269_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT127), .B(G197gat), .Z(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n934_), .A2(new_n630_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n381_), .ZN(G1353gat));
  NOR2_X1   g738(.A1(new_n934_), .A2(new_n673_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AND2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n940_), .B2(new_n941_), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n934_), .B2(new_n666_), .ZN(new_n945_));
  OR2_X1    g744(.A1(new_n662_), .A2(G218gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n934_), .B2(new_n946_), .ZN(G1355gat));
endmodule


