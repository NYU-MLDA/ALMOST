//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT89), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT22), .B1(new_n206_), .B2(KEYINPUT88), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n206_), .A2(KEYINPUT22), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n207_), .B(new_n210_), .C1(new_n211_), .C2(KEYINPUT88), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n205_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n204_), .A2(KEYINPUT89), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT87), .B1(new_n203_), .B2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n203_), .A2(KEYINPUT87), .A3(new_n217_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n208_), .A2(new_n215_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(G190gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n222_), .B(new_n225_), .C1(new_n226_), .C2(new_n223_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n221_), .A3(new_n227_), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n213_), .A2(new_n214_), .B1(new_n218_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G227gat), .A2(G233gat), .ZN(new_n233_));
  INV_X1    g032(.A(G15gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n232_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT31), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT90), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT91), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n238_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n238_), .B(new_n245_), .C1(KEYINPUT91), .C2(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G155gat), .B(G162gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT92), .ZN(new_n250_));
  INV_X1    g049(.A(G141gat), .ZN(new_n251_));
  INV_X1    g050(.A(G148gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT3), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(KEYINPUT3), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n254_), .A2(new_n257_), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n250_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G155gat), .ZN(new_n262_));
  INV_X1    g061(.A(G162gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT1), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(G155gat), .B2(G162gat), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT1), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n255_), .B(new_n253_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n261_), .A2(KEYINPUT93), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT93), .B1(new_n261_), .B2(new_n267_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT29), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n273_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G22gat), .B(G50gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G197gat), .B(G204gat), .Z(new_n282_));
  INV_X1    g081(.A(KEYINPUT94), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT21), .ZN(new_n284_));
  XOR2_X1   g083(.A(G211gat), .B(G218gat), .Z(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n269_), .A2(new_n271_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n289_), .B(new_n290_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n289_), .B(KEYINPUT95), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n261_), .A2(new_n267_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(new_n292_), .ZN(new_n296_));
  OAI211_X1 g095(.A(G228gat), .B(G233gat), .C1(new_n294_), .C2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G78gat), .B(G106gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT96), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n298_), .B(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n281_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n281_), .A2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT101), .ZN(new_n306_));
  INV_X1    g105(.A(new_n241_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n269_), .A2(new_n306_), .A3(new_n271_), .A4(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n268_), .A2(new_n270_), .A3(new_n241_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n295_), .A2(new_n241_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT101), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n291_), .A2(KEYINPUT4), .A3(new_n241_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n312_), .B2(KEYINPUT4), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n317_), .B2(new_n313_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G1gat), .B(G29gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G85gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT0), .B(G57gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n313_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n323_), .A2(KEYINPUT33), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT19), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT22), .B(G169gat), .Z(new_n334_));
  OAI211_X1 g133(.A(new_n204_), .B(new_n209_), .C1(G176gat), .C2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n336_));
  OR3_X1    g135(.A1(new_n336_), .A2(G169gat), .A3(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n220_), .A2(new_n336_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n226_), .A2(new_n222_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n203_), .A4(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n289_), .A2(new_n341_), .A3(KEYINPUT99), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT99), .B1(new_n289_), .B2(new_n341_), .ZN(new_n343_));
  AOI211_X1 g142(.A(new_n331_), .B(new_n333_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n229_), .A2(new_n289_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT98), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT100), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n347_), .A3(KEYINPUT100), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n331_), .B1(new_n289_), .B2(new_n341_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(new_n289_), .B2(new_n229_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n354_), .A2(new_n333_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n330_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n330_), .ZN(new_n358_));
  AOI211_X1 g157(.A(new_n355_), .B(new_n358_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n326_), .B(new_n360_), .C1(KEYINPUT33), .C2(new_n323_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n318_), .A2(new_n322_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n318_), .A2(new_n322_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n354_), .A2(new_n333_), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT102), .Z(new_n367_));
  INV_X1    g166(.A(new_n333_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n341_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n331_), .B1(new_n294_), .B2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n347_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n365_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n352_), .A2(new_n356_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n364_), .B(new_n372_), .C1(new_n373_), .C2(new_n365_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n305_), .B1(new_n361_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n358_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n378_), .B(KEYINPUT27), .C1(new_n373_), .C2(new_n358_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n305_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n364_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n248_), .B1(new_n375_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n380_), .A2(new_n305_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n248_), .A2(new_n364_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G99gat), .A2(G106gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT65), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT6), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT65), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(KEYINPUT65), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(KEYINPUT6), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(G99gat), .A4(G106gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT66), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT7), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G99gat), .A2(G106gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(KEYINPUT67), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT67), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n403_), .A2(G99gat), .A3(G106gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT68), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(KEYINPUT67), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n403_), .B1(G99gat), .B2(G106gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT68), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .A4(new_n400_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n393_), .A2(KEYINPUT66), .A3(new_n396_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n399_), .A2(new_n410_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G85gat), .B(G92gat), .Z(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT8), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n405_), .A2(new_n409_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n393_), .A2(new_n396_), .A3(new_n412_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT69), .B(new_n414_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT8), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n393_), .A2(new_n396_), .A3(new_n412_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n415_), .B1(new_n422_), .B2(new_n410_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(KEYINPUT69), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n417_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G57gat), .B(G64gat), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n426_), .A2(KEYINPUT11), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(KEYINPUT11), .ZN(new_n428_));
  XOR2_X1   g227(.A(G71gat), .B(G78gat), .Z(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n428_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT10), .B(G99gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT64), .ZN(new_n434_));
  INV_X1    g233(.A(G106gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G85gat), .ZN(new_n437_));
  INV_X1    g236(.A(G92gat), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT9), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n414_), .B2(KEYINPUT9), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(new_n411_), .A3(new_n399_), .A4(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n425_), .A2(new_n432_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(G230gat), .ZN(new_n443_));
  INV_X1    g242(.A(G233gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n441_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n419_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n415_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(KEYINPUT8), .A3(new_n420_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n452_), .B2(new_n417_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT12), .B1(new_n453_), .B2(new_n432_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n455_));
  INV_X1    g254(.A(new_n432_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n423_), .B2(KEYINPUT69), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n458_), .A2(new_n451_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n455_), .B(new_n456_), .C1(new_n459_), .C2(new_n448_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n447_), .B1(new_n454_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n425_), .A2(new_n441_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n456_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n446_), .B1(new_n463_), .B2(new_n442_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G120gat), .B(G148gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT5), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G176gat), .B(G204gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(KEYINPUT70), .B2(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G1gat), .A2(G8gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT14), .ZN(new_n484_));
  INV_X1    g283(.A(G22gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n234_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(G15gat), .A2(G22gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n484_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT81), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n488_), .A2(KEYINPUT81), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n483_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G1gat), .A2(G8gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n495_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n482_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(new_n498_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(KEYINPUT84), .A3(new_n502_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n481_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n501_), .B(KEYINPUT15), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n506_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n502_), .A3(new_n481_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT85), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n511_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n514_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(new_n510_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n480_), .A2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n387_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n453_), .A2(new_n501_), .B1(new_n527_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n462_), .A2(KEYINPUT72), .A3(new_n512_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT72), .ZN(new_n534_));
  INV_X1    g333(.A(new_n512_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n453_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(KEYINPUT35), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n512_), .B1(new_n459_), .B2(new_n448_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n425_), .A2(new_n441_), .A3(new_n501_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n531_), .A2(new_n527_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n538_), .B(KEYINPUT76), .Z(new_n544_));
  NAND4_X1  g343(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT77), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n532_), .A2(new_n547_), .A3(new_n541_), .A4(new_n544_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT79), .ZN(new_n550_));
  XOR2_X1   g349(.A(G190gat), .B(G218gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT73), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT36), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n550_), .B1(new_n549_), .B2(new_n555_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT80), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n554_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT74), .B(KEYINPUT75), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n540_), .A2(new_n546_), .A3(new_n548_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT78), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n546_), .A2(new_n548_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n540_), .A4(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .A4(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n549_), .A2(new_n555_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT79), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n571_), .A2(new_n574_), .A3(new_n561_), .A4(new_n556_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT80), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n561_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT82), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n432_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n506_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT17), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n587_), .B(KEYINPUT17), .Z(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n582_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n578_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n526_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n364_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n594_), .A2(G1gat), .A3(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT38), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n559_), .A2(new_n571_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n480_), .A2(new_n592_), .A3(new_n524_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n595_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n597_), .A2(new_n598_), .A3(new_n605_), .ZN(G1324gat));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n380_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609_));
  AND4_X1   g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .A4(G8gat), .ZN(new_n610_));
  INV_X1    g409(.A(G8gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n608_), .A2(new_n612_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n380_), .A2(new_n611_), .ZN(new_n614_));
  OAI22_X1  g413(.A1(new_n610_), .A2(new_n613_), .B1(new_n594_), .B2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g415(.A(new_n248_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n234_), .B1(new_n603_), .B2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT41), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n234_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n594_), .B2(new_n620_), .ZN(G1326gat));
  XNOR2_X1  g420(.A(new_n305_), .B(KEYINPUT104), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n603_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G22gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT42), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n526_), .A2(new_n485_), .A3(new_n593_), .A4(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1327gat));
  NOR2_X1   g429(.A1(new_n599_), .A2(new_n591_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n526_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(G29gat), .B1(new_n632_), .B2(new_n364_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n387_), .A2(new_n578_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n578_), .B2(KEYINPUT106), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n387_), .B(new_n578_), .C1(KEYINPUT106), .C2(new_n635_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n525_), .A2(new_n592_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT44), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  AOI211_X1 g442(.A(new_n643_), .B(new_n640_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n364_), .A2(G29gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n633_), .B1(new_n645_), .B2(new_n646_), .ZN(G1328gat));
  INV_X1    g446(.A(G36gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n632_), .A2(new_n648_), .A3(new_n380_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT45), .ZN(new_n650_));
  INV_X1    g449(.A(new_n380_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n642_), .A2(new_n644_), .A3(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n648_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n650_), .B(KEYINPUT46), .C1(new_n652_), .C2(new_n648_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1329gat));
  AOI21_X1  g456(.A(G43gat), .B1(new_n632_), .B2(new_n617_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n248_), .A2(new_n236_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n645_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT47), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n632_), .B2(new_n623_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n305_), .A2(G50gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n645_), .B2(new_n664_), .ZN(G1331gat));
  NOR3_X1   g464(.A1(new_n479_), .A2(new_n592_), .A3(new_n523_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n601_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G57gat), .B1(new_n668_), .B2(new_n595_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n479_), .A2(new_n523_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n387_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n593_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n595_), .A2(G57gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(G1332gat));
  OAI21_X1  g473(.A(G64gat), .B1(new_n668_), .B2(new_n651_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT107), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n677_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n672_), .A2(G64gat), .A3(new_n651_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(G1333gat));
  INV_X1    g480(.A(G71gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n667_), .B2(new_n617_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n617_), .A2(new_n682_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n672_), .B2(new_n686_), .ZN(G1334gat));
  INV_X1    g486(.A(G78gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n667_), .B2(new_n623_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT50), .Z(new_n690_));
  NAND2_X1  g489(.A1(new_n623_), .A2(new_n688_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n672_), .B2(new_n691_), .ZN(G1335gat));
  NAND2_X1  g491(.A1(new_n671_), .A2(new_n631_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n437_), .B1(new_n693_), .B2(new_n595_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT109), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n670_), .A2(new_n592_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT110), .Z(new_n697_));
  AND2_X1   g496(.A1(new_n639_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n364_), .A2(G85gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT111), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n695_), .B1(new_n698_), .B2(new_n700_), .ZN(G1336gat));
  INV_X1    g500(.A(new_n693_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n438_), .A3(new_n380_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n698_), .A2(new_n380_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n438_), .ZN(G1337gat));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n434_), .A3(new_n617_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n698_), .A2(new_n617_), .ZN(new_n707_));
  INV_X1    g506(.A(G99gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g509(.A1(new_n702_), .A2(new_n435_), .A3(new_n305_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n639_), .A2(new_n305_), .A3(new_n697_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT52), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(G106gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n712_), .B2(G106gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g516(.A1(new_n505_), .A2(new_n509_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n481_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n503_), .A2(new_n481_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n519_), .B1(new_n720_), .B2(new_n513_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n520_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n461_), .B2(KEYINPUT55), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n445_), .B1(new_n453_), .B2(new_n432_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n455_), .B1(new_n462_), .B2(new_n456_), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT12), .B(new_n432_), .C1(new_n425_), .C2(new_n441_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(KEYINPUT114), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n726_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n454_), .A2(new_n460_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT115), .B1(new_n734_), .B2(new_n442_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n459_), .A2(new_n456_), .A3(new_n448_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n736_), .B(new_n737_), .C1(new_n454_), .C2(new_n460_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n445_), .B1(new_n735_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n461_), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n733_), .A2(new_n739_), .A3(new_n741_), .A4(new_n742_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n743_), .A2(KEYINPUT56), .A3(new_n469_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT56), .B1(new_n743_), .B2(new_n469_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n724_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT118), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(KEYINPUT58), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  OAI221_X1 g548(.A(new_n724_), .B1(new_n747_), .B2(KEYINPUT58), .C1(new_n744_), .C2(new_n745_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n578_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n523_), .A2(new_n471_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n523_), .A2(new_n471_), .A3(KEYINPUT113), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n743_), .A2(new_n469_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n743_), .A2(KEYINPUT56), .A3(new_n469_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n474_), .A2(new_n723_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT57), .B(new_n599_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n751_), .A2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n599_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT117), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(KEYINPUT117), .A3(new_n766_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n591_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n575_), .A2(KEYINPUT80), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n575_), .A2(KEYINPUT80), .ZN(new_n772_));
  INV_X1    g571(.A(new_n577_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n523_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n774_), .A2(new_n591_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(KEYINPUT80), .A3(new_n575_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n778_), .A2(new_n591_), .A3(new_n572_), .A4(new_n775_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT119), .B1(new_n770_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n754_), .A2(new_n755_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n762_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n600_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n788_), .B2(KEYINPUT57), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n789_), .A2(new_n769_), .A3(new_n763_), .A4(new_n751_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n592_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  INV_X1    g591(.A(new_n782_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n384_), .A2(new_n364_), .A3(new_n617_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n783_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(G113gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n523_), .ZN(new_n800_));
  XOR2_X1   g599(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n801_));
  NOR2_X1   g600(.A1(new_n788_), .A2(KEYINPUT57), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n592_), .B1(new_n764_), .B2(new_n802_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n795_), .B(new_n801_), .C1(new_n803_), .C2(new_n793_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n524_), .B(new_n804_), .C1(new_n797_), .C2(KEYINPUT59), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n800_), .B1(new_n805_), .B2(new_n799_), .ZN(G1340gat));
  AOI211_X1 g605(.A(new_n479_), .B(new_n804_), .C1(new_n797_), .C2(KEYINPUT59), .ZN(new_n807_));
  INV_X1    g606(.A(G120gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n479_), .B2(KEYINPUT60), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(KEYINPUT60), .B2(new_n808_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n807_), .A2(new_n808_), .B1(new_n797_), .B2(new_n810_), .ZN(G1341gat));
  INV_X1    g610(.A(G127gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n798_), .A2(new_n812_), .A3(new_n591_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n592_), .B(new_n804_), .C1(new_n797_), .C2(KEYINPUT59), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n812_), .ZN(G1342gat));
  AOI21_X1  g614(.A(G134gat), .B1(new_n798_), .B2(new_n600_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n804_), .B1(new_n797_), .B2(KEYINPUT59), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT121), .B(G134gat), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n774_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n816_), .B1(new_n817_), .B2(new_n819_), .ZN(G1343gat));
  NAND2_X1  g619(.A1(new_n783_), .A2(new_n794_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n248_), .A2(new_n305_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n822_), .A2(new_n595_), .A3(new_n380_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n821_), .A2(new_n524_), .A3(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(new_n251_), .ZN(G1344gat));
  NOR3_X1   g625(.A1(new_n821_), .A2(new_n479_), .A3(new_n824_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(new_n252_), .ZN(G1345gat));
  NAND4_X1  g627(.A1(new_n783_), .A2(new_n591_), .A3(new_n794_), .A4(new_n823_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT61), .B(G155gat), .Z(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n792_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n833_));
  AOI211_X1 g632(.A(KEYINPUT119), .B(new_n782_), .C1(new_n790_), .C2(new_n592_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n830_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n835_), .A2(new_n591_), .A3(new_n823_), .A4(new_n836_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n831_), .A2(new_n832_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n831_), .B2(new_n837_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1346gat));
  NAND4_X1  g639(.A1(new_n835_), .A2(new_n263_), .A3(new_n600_), .A4(new_n823_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n821_), .A2(new_n774_), .A3(new_n824_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n263_), .ZN(G1347gat));
  NAND2_X1  g642(.A1(new_n803_), .A2(new_n793_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n385_), .A2(new_n380_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n623_), .A2(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n844_), .A2(new_n523_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n848_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(G169gat), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n334_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n847_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n849_), .A2(KEYINPUT62), .A3(new_n850_), .A4(G169gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(G1348gat));
  AND2_X1   g656(.A1(new_n844_), .A2(new_n846_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G176gat), .B1(new_n858_), .B2(new_n480_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n821_), .A2(new_n305_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n845_), .A2(new_n207_), .A3(new_n479_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1349gat));
  NAND4_X1  g661(.A1(new_n860_), .A2(new_n591_), .A3(new_n380_), .A4(new_n385_), .ZN(new_n863_));
  INV_X1    g662(.A(G183gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n592_), .A2(new_n222_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n863_), .A2(new_n864_), .B1(new_n858_), .B2(new_n865_), .ZN(G1350gat));
  NAND2_X1  g665(.A1(new_n600_), .A2(new_n226_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT125), .Z(new_n868_));
  NAND2_X1  g667(.A1(new_n858_), .A2(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n858_), .A2(new_n578_), .ZN(new_n870_));
  INV_X1    g669(.A(G190gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1351gat));
  NAND3_X1  g671(.A1(new_n248_), .A2(new_n595_), .A3(new_n305_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n651_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n835_), .A2(new_n523_), .A3(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT126), .B(G197gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n835_), .A2(new_n874_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  OAI22_X1  g678(.A1(new_n878_), .A2(new_n479_), .B1(new_n879_), .B2(G204gat), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT127), .B(G204gat), .Z(new_n881_));
  NAND4_X1  g680(.A1(new_n835_), .A2(new_n480_), .A3(new_n874_), .A4(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1353gat));
  NAND3_X1  g682(.A1(new_n835_), .A2(new_n591_), .A3(new_n874_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  AND2_X1   g684(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n884_), .B2(new_n885_), .ZN(G1354gat));
  OAI21_X1  g687(.A(G218gat), .B1(new_n878_), .B2(new_n774_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n599_), .A2(G218gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n878_), .B2(new_n890_), .ZN(G1355gat));
endmodule


