//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n964_, new_n965_,
    new_n967_, new_n968_, new_n969_, new_n971_, new_n972_, new_n973_,
    new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G1gat), .B(G29gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  AND3_X1   g007(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT87), .ZN(new_n213_));
  OAI22_X1  g012(.A1(new_n213_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT87), .B1(new_n215_), .B2(KEYINPUT86), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(KEYINPUT86), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n218_), .A2(new_n213_), .A3(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n211_), .B(new_n212_), .C1(new_n217_), .C2(new_n220_), .ZN(new_n221_));
  OR3_X1    g020(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT85), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n224_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n228_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT1), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(new_n234_), .A3(new_n228_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n233_), .A2(new_n222_), .A3(new_n235_), .A4(new_n223_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n209_), .A2(new_n210_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(new_n219_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n230_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n221_), .A2(new_n229_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT98), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(KEYINPUT98), .A3(new_n244_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n248_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n252_), .A3(KEYINPUT4), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT99), .ZN(new_n255_));
  OR3_X1    g054(.A1(new_n248_), .A2(KEYINPUT4), .A3(new_n245_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n255_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n247_), .A2(new_n252_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n207_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT104), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n207_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT104), .B1(new_n266_), .B2(new_n257_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n261_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT97), .ZN(new_n269_));
  OR2_X1    g068(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(G197gat), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(G204gat), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT92), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n272_), .A2(new_n275_), .A3(KEYINPUT92), .A4(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n273_), .A2(new_n274_), .ZN(new_n284_));
  INV_X1    g083(.A(G204gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT91), .B(G204gat), .ZN(new_n287_));
  INV_X1    g086(.A(G197gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n283_), .B1(new_n290_), .B2(KEYINPUT21), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n281_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n272_), .A2(new_n275_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n282_), .A2(new_n276_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  INV_X1    g100(.A(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n300_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G169gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT22), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n310_), .A2(KEYINPUT96), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT96), .B1(new_n310_), .B2(new_n311_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n304_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n305_), .A2(new_n309_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(KEYINPUT24), .A3(new_n311_), .ZN(new_n319_));
  OR3_X1    g118(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G183gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n302_), .A2(KEYINPUT26), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n327_));
  AND4_X1   g126(.A1(new_n323_), .A2(new_n324_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT95), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT95), .B1(new_n332_), .B2(new_n328_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n314_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n269_), .B1(new_n296_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n295_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n281_), .B2(new_n291_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n304_), .A2(new_n311_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n310_), .A2(KEYINPUT80), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT22), .B(G169gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n309_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n322_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT25), .ZN(new_n346_));
  AND4_X1   g145(.A1(new_n344_), .A2(new_n346_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n332_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n337_), .A2(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n314_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n337_), .A3(KEYINPUT97), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n335_), .A2(new_n350_), .A3(new_n352_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n337_), .A2(new_n349_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n351_), .B2(new_n337_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n354_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G64gat), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(G92gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(G92gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT32), .A3(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n357_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n268_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n321_), .A2(new_n329_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n337_), .A2(new_n370_), .A3(new_n314_), .ZN(new_n371_));
  XOR2_X1   g170(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n337_), .B2(new_n349_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n354_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n355_), .B1(new_n296_), .B2(new_n334_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n354_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n358_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n367_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT103), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n202_), .B1(new_n369_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT103), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n378_), .B(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(KEYINPUT105), .A3(new_n268_), .A4(new_n368_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT94), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT89), .B(G233gat), .Z(new_n387_));
  AND2_X1   g186(.A1(new_n387_), .A2(G228gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT93), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G22gat), .B(G50gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n248_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n248_), .B2(new_n394_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n393_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n397_), .A3(new_n392_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n248_), .A2(new_n394_), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n403_), .A2(new_n337_), .B1(new_n389_), .B2(new_n388_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n386_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n402_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n385_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n365_), .A2(new_n366_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n351_), .A2(KEYINPUT97), .A3(new_n337_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT97), .B1(new_n351_), .B2(new_n337_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n356_), .B1(new_n337_), .B2(new_n349_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n376_), .B1(new_n375_), .B2(new_n358_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n414_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n414_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n357_), .A2(new_n361_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT33), .B1(new_n262_), .B2(new_n264_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n266_), .A2(new_n426_), .A3(new_n257_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n256_), .A2(new_n258_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n207_), .B1(new_n428_), .B2(new_n253_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n247_), .A2(new_n252_), .A3(KEYINPUT101), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT101), .B1(new_n247_), .B2(new_n252_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n255_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n425_), .A2(new_n427_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n413_), .B1(new_n424_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n380_), .A2(new_n383_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n268_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n422_), .A2(KEYINPUT27), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n421_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT27), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT106), .B1(new_n423_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT106), .ZN(new_n443_));
  AOI211_X1 g242(.A(new_n443_), .B(KEYINPUT27), .C1(new_n420_), .C2(new_n422_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n436_), .B(new_n440_), .C1(new_n442_), .C2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n413_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n343_), .B2(new_n348_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n341_), .B1(new_n340_), .B2(new_n309_), .ZN(new_n450_));
  AND4_X1   g249(.A1(new_n341_), .A2(new_n306_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n311_), .B(new_n304_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT26), .B(G190gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n454_), .A2(new_n319_), .A3(new_n317_), .A4(new_n320_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(KEYINPUT30), .A3(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n449_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n449_), .B2(new_n456_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n447_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT81), .Z(new_n463_));
  NOR3_X1   g262(.A1(new_n343_), .A2(new_n348_), .A3(new_n448_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT30), .B1(new_n452_), .B2(new_n455_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n457_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n447_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n449_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n461_), .A2(new_n463_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n463_), .B1(new_n461_), .B2(new_n469_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT31), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n461_), .A2(new_n469_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n463_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT31), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n477_), .A2(new_n471_), .A3(new_n478_), .A4(new_n470_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n245_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n474_), .A2(new_n479_), .A3(new_n246_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n435_), .A2(new_n446_), .A3(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n407_), .A2(new_n412_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n440_), .B(new_n485_), .C1(new_n442_), .C2(new_n444_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n474_), .A2(new_n246_), .A3(new_n479_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n246_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n268_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT107), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n481_), .A2(new_n436_), .A3(new_n482_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT107), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n492_), .A2(new_n486_), .A3(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n484_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT6), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  OR3_X1    g299(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G85gat), .B(G92gat), .Z(new_n503_));
  AOI21_X1  g302(.A(new_n497_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT10), .B(G99gat), .Z(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n499_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT9), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT64), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n503_), .B2(new_n513_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n505_), .A2(new_n506_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  XOR2_X1   g316(.A(G71gat), .B(G78gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(KEYINPUT11), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n511_), .A2(new_n515_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n506_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n525_), .B1(new_n526_), .B2(new_n504_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT65), .B1(new_n527_), .B2(new_n522_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n522_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n529_), .A2(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n527_), .B2(new_n522_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n534_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n285_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT5), .B(G176gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  NAND3_X1  g341(.A1(new_n533_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n496_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n533_), .A2(new_n538_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n542_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT13), .A3(new_n543_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n546_), .A2(new_n550_), .A3(KEYINPUT66), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT66), .B1(new_n546_), .B2(new_n550_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G15gat), .B(G22gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT70), .B(G1gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G8gat), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n557_), .B2(KEYINPUT14), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G1gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(G8gat), .ZN(new_n560_));
  INV_X1    g359(.A(G1gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n558_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(G8gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G29gat), .B(G36gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G43gat), .B(G50gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT74), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT75), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT76), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n569_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT76), .B1(new_n575_), .B2(KEYINPUT75), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n565_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n569_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n574_), .A2(new_n576_), .A3(new_n578_), .A4(new_n569_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n568_), .B(KEYINPUT15), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n578_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n581_), .A3(new_n571_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT78), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT77), .B(G113gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n584_), .A2(new_n587_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n554_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n495_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n601_));
  INV_X1    g400(.A(G231gat), .ZN(new_n602_));
  INV_X1    g401(.A(G233gat), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n560_), .A2(new_n564_), .A3(new_n605_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n522_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n608_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n523_), .B1(new_n610_), .B2(new_n606_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT71), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n609_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(new_n301_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(G211gat), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT17), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n612_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT72), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n609_), .A2(new_n611_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT71), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT72), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n619_), .A4(new_n613_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n617_), .B(new_n618_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n601_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT73), .B(new_n629_), .C1(new_n622_), .C2(new_n626_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n516_), .A2(new_n568_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n527_), .A2(new_n585_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT68), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT67), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT34), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT35), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n644_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n648_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n642_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n641_), .A2(new_n644_), .A3(new_n649_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n638_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n636_), .A2(new_n637_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n652_), .A2(new_n637_), .A3(new_n636_), .A4(new_n653_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(KEYINPUT69), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT37), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n600_), .A2(new_n633_), .A3(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n436_), .A2(new_n556_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT108), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT38), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n656_), .A2(new_n657_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n495_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n627_), .A2(new_n630_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n554_), .A2(new_n598_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G1gat), .B1(new_n669_), .B2(new_n436_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n664_), .A2(new_n670_), .ZN(G1324gat));
  NOR3_X1   g470(.A1(new_n418_), .A2(new_n419_), .A3(new_n414_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n421_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n441_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n443_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n423_), .A2(KEYINPUT106), .A3(new_n441_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n439_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n660_), .A2(new_n563_), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G8gat), .B1(new_n669_), .B2(new_n677_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT39), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT39), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n483_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n660_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT109), .Z(new_n688_));
  OAI21_X1  g487(.A(G15gat), .B1(new_n669_), .B2(new_n483_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT41), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(KEYINPUT41), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n690_), .A3(new_n691_), .ZN(G1326gat));
  OAI21_X1  g491(.A(G22gat), .B1(new_n669_), .B2(new_n485_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT42), .ZN(new_n694_));
  INV_X1    g493(.A(G22gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n660_), .A2(new_n695_), .A3(new_n413_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n633_), .A2(new_n665_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n600_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(G29gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n268_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n633_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n599_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n659_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n495_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT43), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n495_), .A2(new_n707_), .A3(new_n704_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT44), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n713_));
  AOI211_X1 g512(.A(KEYINPUT110), .B(new_n703_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n268_), .B(new_n710_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G29gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n715_), .A2(new_n716_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n701_), .B1(new_n718_), .B2(new_n719_), .ZN(G1328gat));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT114), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT115), .Z(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n677_), .A2(G36gat), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n698_), .A2(new_n495_), .A3(new_n599_), .A4(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n727_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n728_), .A2(new_n731_), .A3(new_n729_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n677_), .B1(new_n709_), .B2(KEYINPUT44), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n737_), .B2(G36gat), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n721_), .A2(KEYINPUT114), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n724_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n739_), .ZN(new_n741_));
  INV_X1    g540(.A(G36gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n706_), .A2(new_n708_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n703_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT110), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n709_), .A2(new_n712_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n711_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n742_), .B1(new_n748_), .B2(new_n736_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n741_), .B(new_n723_), .C1(new_n749_), .C2(new_n735_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n740_), .A2(new_n750_), .ZN(G1329gat));
  NAND4_X1  g550(.A1(new_n748_), .A2(G43gat), .A3(new_n686_), .A4(new_n710_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n699_), .A2(new_n686_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(G43gat), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n752_), .A2(new_n757_), .A3(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1330gat));
  AOI21_X1  g558(.A(G50gat), .B1(new_n699_), .B2(new_n413_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n748_), .A2(new_n710_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n413_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1331gat));
  OAI211_X1 g562(.A(new_n594_), .B(new_n596_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n495_), .A2(new_n633_), .A3(new_n659_), .A4(new_n765_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n766_), .A2(G57gat), .A3(new_n436_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n764_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n495_), .A2(new_n665_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT116), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n495_), .A2(new_n768_), .A3(new_n771_), .A4(new_n665_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n268_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n767_), .B1(new_n774_), .B2(G57gat), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT117), .ZN(G1332gat));
  OR3_X1    g575(.A1(new_n766_), .A2(G64gat), .A3(new_n677_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n678_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G64gat), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT48), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT48), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1333gat));
  OR3_X1    g581(.A1(new_n766_), .A2(G71gat), .A3(new_n483_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n686_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G71gat), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(KEYINPUT49), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(KEYINPUT49), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1334gat));
  OR3_X1    g587(.A1(new_n766_), .A2(G78gat), .A3(new_n485_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n770_), .A2(new_n413_), .A3(new_n772_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(G78gat), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n790_), .B2(G78gat), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n790_), .A2(G78gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT118), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT50), .B1(new_n798_), .B2(new_n792_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n789_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT119), .B(new_n789_), .C1(new_n796_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1335gat));
  NOR3_X1   g603(.A1(new_n633_), .A2(new_n665_), .A3(new_n764_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n495_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G85gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n268_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n633_), .B(new_n764_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(new_n268_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(new_n808_), .ZN(G1336gat));
  INV_X1    g611(.A(G92gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n807_), .A2(new_n813_), .A3(new_n678_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n810_), .A2(new_n678_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n813_), .ZN(G1337gat));
  AND2_X1   g615(.A1(new_n810_), .A2(new_n686_), .ZN(new_n817_));
  INV_X1    g616(.A(G99gat), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n686_), .A2(new_n507_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n817_), .A2(new_n818_), .B1(new_n806_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g620(.A1(new_n807_), .A2(new_n508_), .A3(new_n413_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n810_), .A2(new_n413_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(G106gat), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT52), .B(new_n508_), .C1(new_n810_), .C2(new_n413_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n822_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT53), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n829_), .B(new_n822_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1339gat));
  NOR3_X1   g630(.A1(new_n483_), .A2(new_n486_), .A3(new_n436_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n667_), .A2(KEYINPUT73), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n584_), .A2(new_n587_), .A3(new_n595_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n595_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n546_), .A2(new_n550_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n627_), .A2(new_n601_), .A3(new_n630_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n834_), .A2(new_n659_), .A3(new_n838_), .A4(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT120), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n633_), .A2(new_n842_), .A3(new_n659_), .A4(new_n838_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n841_), .A2(KEYINPUT54), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT54), .B1(new_n841_), .B2(new_n843_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n528_), .B(new_n524_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n847_), .A2(new_n532_), .B1(new_n538_), .B2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT55), .B(new_n534_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n542_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT122), .B1(new_n851_), .B2(KEYINPUT56), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n532_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n538_), .A2(new_n848_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n850_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n548_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n852_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n851_), .A2(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n580_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n575_), .A2(new_n581_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n595_), .B1(new_n864_), .B2(new_n586_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n596_), .A2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n862_), .A2(KEYINPUT58), .A3(new_n543_), .A4(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n852_), .A2(new_n859_), .B1(KEYINPUT56), .B2(new_n851_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n596_), .A2(new_n543_), .A3(new_n866_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n868_), .A2(new_n872_), .A3(new_n704_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n665_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n856_), .A2(new_n858_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n544_), .B1(new_n861_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n549_), .A2(new_n543_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n596_), .A2(new_n877_), .A3(new_n866_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n597_), .A2(new_n876_), .B1(new_n878_), .B2(KEYINPUT121), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n878_), .A2(KEYINPUT121), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n874_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n873_), .B1(new_n881_), .B2(KEYINPUT57), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n883_), .B(new_n874_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n667_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n833_), .B1(new_n846_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT59), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n702_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n846_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n832_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G113gat), .B1(new_n893_), .B2(new_n598_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n886_), .B(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n598_), .A2(G113gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n894_), .B1(new_n897_), .B2(new_n898_), .ZN(G1340gat));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n553_), .B2(G120gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n892_), .B(new_n554_), .C1(new_n891_), .C2(new_n886_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n896_), .B2(new_n901_), .ZN(new_n904_));
  INV_X1    g703(.A(G120gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n904_), .B2(new_n905_), .ZN(G1341gat));
  OAI21_X1  g705(.A(G127gat), .B1(new_n893_), .B2(new_n667_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n702_), .A2(G127gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n897_), .B2(new_n908_), .ZN(G1342gat));
  NAND2_X1  g708(.A1(new_n896_), .A2(new_n874_), .ZN(new_n910_));
  INV_X1    g709(.A(G134gat), .ZN(new_n911_));
  INV_X1    g710(.A(new_n893_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n704_), .A2(G134gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT124), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n910_), .A2(new_n911_), .B1(new_n912_), .B2(new_n914_), .ZN(G1343gat));
  NAND2_X1  g714(.A1(new_n846_), .A2(new_n885_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n686_), .A2(new_n678_), .A3(new_n436_), .A4(new_n485_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(KEYINPUT125), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(KEYINPUT125), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n597_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(G141gat), .ZN(new_n922_));
  INV_X1    g721(.A(G141gat), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n923_), .B(new_n597_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1344gat));
  OAI21_X1  g724(.A(new_n554_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G148gat), .ZN(new_n927_));
  INV_X1    g726(.A(G148gat), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n928_), .B(new_n554_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1345gat));
  OAI21_X1  g729(.A(new_n633_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT61), .B(G155gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n932_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n633_), .B(new_n934_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1346gat));
  INV_X1    g735(.A(new_n920_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n918_), .A2(KEYINPUT125), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n659_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(G162gat), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n919_), .A2(new_n920_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n874_), .A2(new_n940_), .ZN(new_n942_));
  OAI22_X1  g741(.A1(new_n939_), .A2(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1347gat));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n678_), .A2(new_n490_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n413_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n846_), .B2(new_n889_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n948_), .A2(new_n597_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n944_), .B1(new_n949_), .B2(new_n305_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n305_), .B1(new_n948_), .B2(new_n597_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(KEYINPUT62), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n948_), .A2(new_n340_), .A3(new_n597_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n950_), .A2(new_n951_), .A3(new_n953_), .A4(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n952_), .B2(KEYINPUT62), .ZN(new_n956_));
  AOI211_X1 g755(.A(new_n944_), .B(new_n305_), .C1(new_n948_), .C2(new_n597_), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT126), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n955_), .A2(new_n958_), .ZN(G1348gat));
  AOI21_X1  g758(.A(G176gat), .B1(new_n948_), .B2(new_n554_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n413_), .B1(new_n846_), .B2(new_n885_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n945_), .A2(new_n553_), .A3(new_n309_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n960_), .B1(new_n961_), .B2(new_n962_), .ZN(G1349gat));
  NAND4_X1  g762(.A1(new_n961_), .A2(new_n678_), .A3(new_n490_), .A4(new_n633_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n667_), .B1(new_n323_), .B2(new_n327_), .ZN(new_n965_));
  AOI22_X1  g764(.A1(new_n964_), .A2(new_n301_), .B1(new_n948_), .B2(new_n965_), .ZN(G1350gat));
  INV_X1    g765(.A(new_n948_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G190gat), .B1(new_n967_), .B2(new_n659_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n948_), .A2(new_n874_), .A3(new_n453_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1351gat));
  NAND3_X1  g769(.A1(new_n678_), .A2(new_n436_), .A3(new_n413_), .ZN(new_n971_));
  AOI211_X1 g770(.A(new_n686_), .B(new_n971_), .C1(new_n846_), .C2(new_n885_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(new_n597_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g773(.A1(new_n972_), .A2(new_n554_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n975_), .A2(G204gat), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n976_), .B1(new_n287_), .B2(new_n975_), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n972_), .A2(new_n627_), .A3(new_n630_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n979_));
  AND2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n978_), .A2(new_n979_), .A3(new_n980_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n978_), .B2(new_n979_), .ZN(G1354gat));
  INV_X1    g781(.A(G218gat), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n972_), .A2(new_n983_), .A3(new_n874_), .ZN(new_n984_));
  AND2_X1   g783(.A1(new_n972_), .A2(new_n704_), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n984_), .B1(new_n985_), .B2(new_n983_), .ZN(G1355gat));
endmodule


