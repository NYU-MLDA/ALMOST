//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_;
  XNOR2_X1  g000(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n202_));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203_));
  INV_X1    g002(.A(G155gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT1), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G155gat), .B2(G162gat), .ZN(new_n207_));
  NOR3_X1   g006(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT1), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n203_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT84), .ZN(new_n210_));
  NOR3_X1   g009(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT85), .Z(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT86), .ZN(new_n214_));
  INV_X1    g013(.A(G141gat), .ZN(new_n215_));
  INV_X1    g014(.A(G148gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n217_), .A2(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(KEYINPUT2), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n212_), .A2(new_n214_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT87), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n224_), .A3(new_n221_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n210_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G22gat), .B(G50gat), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n202_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n232_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n202_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n230_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G197gat), .B(G204gat), .Z(new_n238_));
  XOR2_X1   g037(.A(G211gat), .B(G218gat), .Z(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT21), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT90), .Z(new_n241_));
  NOR2_X1   g040(.A1(new_n238_), .A2(KEYINPUT21), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(new_n239_), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n245_));
  OAI211_X1 g044(.A(KEYINPUT21), .B(new_n245_), .C1(new_n238_), .C2(KEYINPUT89), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G78gat), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n241_), .A2(new_n247_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n210_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n220_), .A2(new_n224_), .A3(new_n221_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n224_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(KEYINPUT29), .ZN(new_n256_));
  INV_X1    g055(.A(G78gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(new_n258_), .A3(G106gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(G106gat), .B1(new_n250_), .B2(new_n258_), .ZN(new_n261_));
  OAI211_X1 g060(.A(G228gat), .B(G233gat), .C1(new_n251_), .C2(KEYINPUT91), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n250_), .A2(new_n258_), .ZN(new_n265_));
  INV_X1    g064(.A(G106gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n262_), .B1(new_n267_), .B2(new_n259_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n237_), .B1(new_n264_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n237_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n263_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT78), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT24), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT78), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n276_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT24), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT23), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT25), .B(G183gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT77), .B(G190gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT26), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n287_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n284_), .A2(new_n286_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT79), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(KEYINPUT22), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT22), .B(G169gat), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n294_), .B(new_n297_), .C1(new_n298_), .C2(new_n295_), .ZN(new_n299_));
  INV_X1    g098(.A(G183gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n288_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n285_), .B(KEYINPUT23), .Z(new_n302_));
  OAI211_X1 g101(.A(new_n278_), .B(new_n299_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n293_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n275_), .B1(new_n304_), .B2(new_n251_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n287_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n284_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT95), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n302_), .B2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n286_), .B(KEYINPUT95), .C1(G183gat), .C2(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n278_), .A2(KEYINPUT94), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n278_), .A2(KEYINPUT94), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n314_), .A2(new_n315_), .B1(new_n298_), .B2(new_n294_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n248_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT96), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT96), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n248_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n305_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT93), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n304_), .A2(new_n251_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT20), .B1(new_n318_), .B2(new_n248_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n326_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT18), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n328_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT27), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT98), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n329_), .B1(new_n343_), .B2(new_n330_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n330_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT98), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n326_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  OAI22_X1  g146(.A1(new_n347_), .A2(KEYINPUT99), .B1(new_n323_), .B2(new_n327_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n304_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n248_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(new_n345_), .B2(KEYINPUT98), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n330_), .A2(new_n343_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n331_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT99), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n339_), .B1(new_n348_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n341_), .A2(KEYINPUT27), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n342_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT81), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n361_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT82), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT82), .B1(new_n362_), .B2(new_n364_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n360_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n375_), .A2(KEYINPUT83), .A3(new_n371_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n255_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n226_), .A2(new_n369_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT4), .ZN(new_n379_));
  INV_X1    g178(.A(new_n376_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT83), .B1(new_n375_), .B2(new_n371_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n255_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(KEYINPUT97), .Z(new_n386_));
  NAND3_X1  g185(.A1(new_n379_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n377_), .A2(new_n378_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n386_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392_));
  INV_X1    g191(.A(G85gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT0), .B(G57gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n399_), .A2(KEYINPUT100), .A3(new_n387_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT100), .B1(new_n399_), .B2(new_n387_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n349_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n349_), .A2(new_n406_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(new_n382_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(KEYINPUT80), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT30), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT31), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n410_), .B(new_n414_), .ZN(new_n415_));
  AND4_X1   g214(.A1(new_n274_), .A2(new_n359_), .A3(new_n403_), .A4(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT32), .B(new_n338_), .C1(new_n348_), .C2(new_n355_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n338_), .A2(KEYINPUT32), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n328_), .A2(new_n333_), .A3(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n402_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT101), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT101), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n402_), .A2(new_n417_), .A3(new_n422_), .A4(new_n419_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n340_), .A2(new_n341_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n377_), .A2(new_n378_), .A3(new_n386_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n397_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n384_), .A2(new_n389_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n379_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n399_), .A2(KEYINPUT33), .A3(new_n387_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT33), .B1(new_n399_), .B2(new_n387_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n269_), .A2(new_n273_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n421_), .A2(new_n423_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n359_), .A2(new_n403_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n269_), .A2(new_n273_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n415_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n416_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT10), .B(G99gat), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n266_), .ZN(new_n440_));
  INV_X1    g239(.A(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n393_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G85gat), .A2(G92gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT9), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n443_), .A2(KEYINPUT9), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n440_), .A2(new_n444_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n442_), .A2(KEYINPUT64), .A3(new_n443_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI211_X1 g255(.A(KEYINPUT8), .B(new_n452_), .C1(new_n456_), .C2(new_n449_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n266_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n447_), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n453_), .B(new_n461_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n452_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n451_), .B1(new_n457_), .B2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G29gat), .B(G36gat), .Z(new_n468_));
  XOR2_X1   g267(.A(G43gat), .B(G50gat), .Z(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  OR3_X1    g269(.A1(new_n467_), .A2(KEYINPUT66), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT66), .B1(new_n467_), .B2(new_n470_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT35), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G232gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT34), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n471_), .A2(new_n472_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n470_), .B(KEYINPUT15), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n467_), .A2(KEYINPUT65), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n480_), .B(new_n451_), .C1(new_n457_), .C2(new_n466_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n476_), .A2(new_n473_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n484_), .A2(KEYINPUT67), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n477_), .A2(KEYINPUT67), .A3(new_n484_), .A4(new_n482_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G190gat), .B(G218gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G134gat), .B(G162gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT36), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT68), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  AOI211_X1 g299(.A(new_n499_), .B(new_n500_), .C1(new_n491_), .C2(new_n492_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT69), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  AOI211_X1 g301(.A(new_n487_), .B(new_n489_), .C1(new_n477_), .C2(new_n482_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n492_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n497_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n499_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT69), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n493_), .A2(KEYINPUT68), .A3(new_n497_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n496_), .B(KEYINPUT36), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT70), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n491_), .A2(new_n492_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT71), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n502_), .A2(new_n509_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT37), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(new_n512_), .C1(new_n498_), .C2(new_n501_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT72), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n506_), .A2(new_n508_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT72), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n516_), .A4(new_n512_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(KEYINPUT11), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n526_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G1gat), .ZN(new_n534_));
  INV_X1    g333(.A(G8gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT73), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(KEYINPUT73), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G8gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT74), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n542_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n533_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT16), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT17), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n548_), .B(new_n553_), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n546_), .A2(KEYINPUT17), .A3(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT76), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n523_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n478_), .A2(new_n545_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n470_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n545_), .A2(new_n470_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n566_), .B2(new_n562_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G169gat), .B(G197gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n567_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n531_), .B(new_n451_), .C1(new_n457_), .C2(new_n466_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT12), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n529_), .A2(new_n530_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n467_), .A2(new_n526_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(KEYINPUT12), .B(new_n526_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n479_), .A2(new_n481_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n577_), .A2(new_n574_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G120gat), .B(G148gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT5), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n589_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(KEYINPUT13), .A3(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR4_X1   g395(.A1(new_n438_), .A2(new_n558_), .A3(new_n573_), .A4(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n534_), .A3(new_n402_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n519_), .A2(new_n512_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n438_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n556_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n605_), .A2(new_n596_), .A3(new_n573_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n403_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n601_), .A3(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n607_), .B2(new_n359_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n359_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n604_), .A2(KEYINPUT103), .A3(new_n612_), .A4(new_n606_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(G8gat), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT104), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT39), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n611_), .A2(new_n617_), .A3(G8gat), .A4(new_n613_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(KEYINPUT39), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n597_), .A2(new_n535_), .A3(new_n612_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n616_), .A2(KEYINPUT40), .A3(new_n619_), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  INV_X1    g424(.A(new_n415_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G15gat), .B1(new_n607_), .B2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT105), .Z(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n630_));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n597_), .A2(new_n631_), .A3(new_n415_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n630_), .A3(new_n632_), .ZN(G1326gat));
  OAI21_X1  g432(.A(G22gat), .B1(new_n607_), .B2(new_n274_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n597_), .A2(new_n636_), .A3(new_n436_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1327gat));
  INV_X1    g437(.A(new_n557_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n596_), .A2(new_n573_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n639_), .B(new_n640_), .C1(KEYINPUT107), .C2(KEYINPUT44), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n434_), .A2(new_n437_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n416_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n523_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n438_), .A2(KEYINPUT43), .A3(new_n523_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n642_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT107), .B1(KEYINPUT106), .B2(KEYINPUT44), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n646_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT43), .B1(new_n438_), .B2(new_n523_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n642_), .A3(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n402_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n639_), .A2(new_n603_), .ZN(new_n660_));
  NOR4_X1   g459(.A1(new_n438_), .A2(new_n573_), .A3(new_n596_), .A4(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n403_), .A2(G29gat), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n659_), .A2(G29gat), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(G1328gat));
  NAND2_X1  g464(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n666_));
  NOR2_X1   g465(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n668_), .A3(new_n612_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n670_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n651_), .B1(new_n656_), .B2(new_n642_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n641_), .B(new_n652_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n674_), .B(new_n612_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n658_), .B2(new_n612_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n666_), .B(new_n673_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n612_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT109), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(G36gat), .A3(new_n677_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n666_), .B1(new_n684_), .B2(new_n673_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n681_), .A2(new_n685_), .ZN(G1329gat));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n661_), .A2(new_n687_), .A3(new_n415_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n626_), .B1(new_n653_), .B2(new_n657_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n687_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n690_), .B(new_n691_), .Z(G1330gat));
  AOI21_X1  g491(.A(G50gat), .B1(new_n661_), .B2(new_n436_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n436_), .A2(G50gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n658_), .B2(new_n694_), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n438_), .A2(new_n572_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n696_), .A2(new_n596_), .A3(new_n557_), .A4(new_n523_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(G57gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n402_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n596_), .A2(new_n573_), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n438_), .A2(new_n639_), .A3(new_n603_), .A4(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(new_n402_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n703_), .B2(new_n699_), .ZN(G1332gat));
  INV_X1    g503(.A(G64gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n702_), .B2(new_n612_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n698_), .A2(new_n705_), .A3(new_n612_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n702_), .B2(new_n415_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT49), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n698_), .A2(new_n711_), .A3(new_n415_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1334gat));
  AOI21_X1  g514(.A(new_n257_), .B1(new_n702_), .B2(new_n436_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT50), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n698_), .A2(new_n257_), .A3(new_n436_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n557_), .A2(new_n701_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n656_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n403_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n596_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n660_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n696_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n393_), .A3(new_n402_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n728_), .ZN(G1336gat));
  OAI21_X1  g528(.A(G92gat), .B1(new_n722_), .B2(new_n359_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(new_n441_), .A3(new_n612_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n722_), .B2(new_n626_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n415_), .A3(new_n439_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT51), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n735_), .B(new_n737_), .Z(G1338gat));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n266_), .A3(new_n436_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n721_), .A2(new_n436_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G106gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT52), .B(new_n266_), .C1(new_n721_), .C2(new_n436_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g544(.A1(new_n523_), .A2(new_n573_), .A3(new_n724_), .A4(new_n557_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n567_), .A2(new_n571_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n559_), .A2(G229gat), .A3(G233gat), .A4(new_n561_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n570_), .B1(new_n565_), .B2(new_n562_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n582_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(KEYINPUT55), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n583_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT115), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n583_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n589_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n590_), .B(new_n752_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n647_), .A2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n572_), .A2(new_n590_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n764_), .B2(KEYINPUT116), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n770_), .B(KEYINPUT56), .C1(new_n761_), .C2(new_n589_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT117), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n768_), .B(new_n774_), .C1(new_n769_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n752_), .A2(new_n592_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n602_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT57), .B1(new_n778_), .B2(KEYINPUT118), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  AOI211_X1 g580(.A(new_n780_), .B(new_n781_), .C1(new_n777_), .C2(new_n602_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n767_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n748_), .B1(new_n783_), .B2(new_n605_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n436_), .A2(new_n612_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n626_), .A2(new_n403_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT59), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n746_), .B(KEYINPUT54), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n647_), .A2(new_n766_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n772_), .A2(KEYINPUT117), .B1(new_n592_), .B2(new_n752_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n603_), .B1(new_n792_), .B2(new_n775_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n781_), .B1(new_n793_), .B2(new_n780_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n778_), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n790_), .B1(new_n796_), .B2(new_n556_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n787_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(KEYINPUT59), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n789_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n796_), .B2(new_n557_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n783_), .A2(KEYINPUT120), .A3(new_n639_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n790_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n787_), .A2(KEYINPUT59), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT121), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n810_), .A3(new_n807_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n802_), .A2(new_n572_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G113gat), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n799_), .A2(G113gat), .A3(new_n573_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1340gat));
  NAND4_X1  g614(.A1(new_n802_), .A2(new_n596_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G120gat), .ZN(new_n817_));
  INV_X1    g616(.A(new_n799_), .ZN(new_n818_));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n724_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n818_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n819_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(G1341gat));
  NAND4_X1  g621(.A1(new_n802_), .A2(new_n556_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G127gat), .ZN(new_n824_));
  OR3_X1    g623(.A1(new_n799_), .A2(G127gat), .A3(new_n639_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1342gat));
  NAND4_X1  g625(.A1(new_n802_), .A2(new_n647_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G134gat), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n799_), .A2(G134gat), .A3(new_n602_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n436_), .A2(new_n626_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n784_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n359_), .A3(new_n402_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n573_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n215_), .ZN(G1344gat));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n724_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(new_n216_), .ZN(G1345gat));
  NOR2_X1   g636(.A1(new_n833_), .A2(new_n639_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT61), .B(G155gat), .Z(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1346gat));
  OAI21_X1  g639(.A(G162gat), .B1(new_n833_), .B2(new_n523_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n603_), .A2(new_n205_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n833_), .B2(new_n842_), .ZN(G1347gat));
  NOR2_X1   g642(.A1(new_n359_), .A2(new_n402_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n415_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n436_), .A3(new_n573_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n296_), .B1(new_n806_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n847_), .A2(new_n848_), .A3(KEYINPUT62), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n806_), .A2(new_n298_), .A3(new_n846_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n847_), .A2(new_n848_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT62), .B1(new_n847_), .B2(new_n848_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n849_), .B(new_n850_), .C1(new_n851_), .C2(new_n852_), .ZN(G1348gat));
  INV_X1    g652(.A(new_n845_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n806_), .A2(new_n274_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n294_), .B1(new_n855_), .B2(new_n724_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n845_), .A2(new_n724_), .A3(new_n294_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n797_), .A2(new_n274_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n856_), .A2(new_n858_), .A3(KEYINPUT123), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1349gat));
  NOR3_X1   g662(.A1(new_n855_), .A2(new_n287_), .A3(new_n605_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n797_), .A2(new_n274_), .A3(new_n557_), .A4(new_n854_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n300_), .B2(new_n865_), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n855_), .B2(new_n523_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n603_), .A2(new_n306_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n855_), .B2(new_n868_), .ZN(G1351gat));
  NAND2_X1  g668(.A1(new_n832_), .A2(new_n844_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n573_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n244_), .ZN(G1352gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n724_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT124), .B(G204gat), .Z(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n873_), .B2(new_n876_), .ZN(G1353gat));
  NAND2_X1  g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n556_), .A2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT125), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n832_), .A2(new_n844_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT126), .ZN(new_n882_));
  NOR2_X1   g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n832_), .A2(new_n884_), .A3(new_n844_), .A4(new_n880_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n883_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1354gat));
  OAI21_X1  g687(.A(G218gat), .B1(new_n870_), .B2(new_n523_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n602_), .A2(G218gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n870_), .B2(new_n890_), .ZN(G1355gat));
endmodule


