//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT89), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(new_n205_), .B2(new_n204_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n205_), .A2(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT89), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n203_), .A2(KEYINPUT90), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n203_), .A2(KEYINPUT90), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n209_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT3), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT2), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  OR3_X1    g020(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n218_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(new_n216_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(KEYINPUT1), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT85), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n222_), .B(new_n223_), .C1(KEYINPUT1), .C2(new_n221_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n227_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT86), .B(new_n227_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n225_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n215_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(G228gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(G228gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n239_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G78gat), .B(G106gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT91), .Z(new_n247_));
  INV_X1    g046(.A(new_n244_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n215_), .B(new_n248_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n249_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(KEYINPUT92), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n247_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT92), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n250_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G22gat), .B(G50gat), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT28), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n236_), .A2(new_n261_), .A3(new_n237_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n263_), .A2(KEYINPUT87), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n236_), .A2(new_n237_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT28), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n268_), .B2(new_n262_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n260_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT87), .B1(new_n263_), .B2(new_n264_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n266_), .A3(new_n262_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n259_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n258_), .A2(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n253_), .A2(new_n250_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT93), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT82), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G127gat), .B(G134gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT83), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n282_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n288_), .B2(new_n287_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n290_), .A2(new_n292_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n295_));
  AOI21_X1  g094(.A(G176gat), .B1(new_n295_), .B2(KEYINPUT22), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G169gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(G183gat), .A3(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(G183gat), .B2(G190gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n297_), .B1(new_n298_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n300_), .B(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(new_n302_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT25), .B(G183gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G190gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n310_), .B(new_n315_), .C1(KEYINPUT24), .C2(new_n313_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n304_), .B1(new_n307_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G227gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(G15gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT30), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n317_), .B(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT81), .B(G43gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n293_), .A2(new_n294_), .A3(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT94), .ZN(new_n330_));
  INV_X1    g129(.A(new_n215_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n316_), .A2(new_n303_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n314_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G169gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n312_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n307_), .B2(new_n298_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n336_), .B2(KEYINPUT95), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT95), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n335_), .C1(new_n307_), .C2(new_n298_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n331_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT20), .B1(new_n215_), .B2(new_n317_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n330_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(new_n331_), .A3(new_n339_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n329_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n215_), .B2(new_n317_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT27), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n336_), .A2(KEYINPUT95), .ZN(new_n354_));
  INV_X1    g153(.A(new_n332_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n339_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n341_), .B1(new_n356_), .B2(new_n215_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n330_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n331_), .A2(new_n336_), .A3(new_n355_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n350_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n357_), .A2(new_n358_), .B1(new_n360_), .B2(new_n329_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(new_n346_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n353_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n346_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n356_), .A2(new_n215_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n341_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n358_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n364_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT27), .B1(new_n369_), .B2(new_n352_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n281_), .A2(new_n327_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n274_), .A2(new_n277_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT93), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT100), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT27), .ZN(new_n379_));
  INV_X1    g178(.A(new_n352_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n346_), .B1(new_n342_), .B2(new_n351_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n352_), .B(KEYINPUT27), .C1(new_n361_), .C2(new_n346_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT100), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n327_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n376_), .A2(new_n276_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n372_), .A2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G1gat), .B(G29gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(G57gat), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT96), .B1(new_n236_), .B2(new_n287_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n234_), .A2(new_n235_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n224_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n286_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(KEYINPUT96), .A3(new_n286_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n397_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n401_), .A2(KEYINPUT4), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n396_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n395_), .A3(new_n403_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n394_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT99), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n394_), .A3(new_n407_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n388_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n342_), .A2(new_n351_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n361_), .B2(new_n415_), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n404_), .A2(new_n396_), .A3(new_n405_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n402_), .A2(new_n403_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n393_), .B1(new_n419_), .B2(new_n396_), .ZN(new_n420_));
  AOI211_X1 g219(.A(new_n380_), .B(new_n381_), .C1(new_n418_), .C2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n408_), .B1(KEYINPUT98), .B2(KEYINPUT33), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n408_), .A2(KEYINPUT98), .A3(KEYINPUT33), .ZN(new_n424_));
  OAI22_X1  g223(.A1(new_n413_), .A2(new_n417_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n376_), .A2(new_n276_), .A3(new_n327_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n414_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT35), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n431_));
  AND3_X1   g230(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT10), .B(G99gat), .Z(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  AOI211_X1 g233(.A(new_n431_), .B(new_n432_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT65), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT9), .ZN(new_n439_));
  INV_X1    g238(.A(G85gat), .ZN(new_n440_));
  INV_X1    g239(.A(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT64), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT64), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G92gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n440_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n436_), .B(new_n439_), .C1(new_n445_), .C2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT64), .B(G92gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n450_), .B2(new_n440_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n436_), .B1(new_n451_), .B2(new_n439_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n435_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G29gat), .B(G36gat), .Z(new_n454_));
  XOR2_X1   g253(.A(G43gat), .B(G50gat), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G29gat), .B(G36gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G43gat), .B(G50gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468_));
  INV_X1    g267(.A(G99gat), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n434_), .A4(KEYINPUT67), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n432_), .A2(new_n431_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n434_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT67), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n467_), .A2(new_n470_), .A3(new_n471_), .A4(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT68), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n437_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT68), .B1(new_n438_), .B2(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n462_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n475_), .A2(new_n462_), .A3(new_n481_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n453_), .B(new_n461_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n474_), .A2(new_n471_), .A3(new_n470_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n465_), .A2(new_n466_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n481_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT8), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n475_), .A2(new_n462_), .A3(new_n481_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n442_), .A2(new_n444_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n447_), .B1(new_n490_), .B2(G85gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n439_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT65), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n448_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n488_), .A2(new_n489_), .B1(new_n494_), .B2(new_n435_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n456_), .A2(KEYINPUT15), .A3(new_n459_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT15), .B1(new_n456_), .B2(new_n459_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n484_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT72), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT73), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n499_), .B2(KEYINPUT73), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n430_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n488_), .A2(new_n489_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n504_), .A2(new_n461_), .A3(new_n453_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n498_), .B1(new_n504_), .B2(new_n453_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT73), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT72), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT73), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT35), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT34), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n499_), .A2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n503_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n513_), .B1(new_n503_), .B2(new_n510_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G134gat), .B(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT36), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n515_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n519_), .B(KEYINPUT36), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n501_), .A2(new_n502_), .A3(new_n430_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT35), .B1(new_n508_), .B2(new_n509_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n512_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n503_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT37), .B1(new_n522_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT74), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT75), .B1(new_n515_), .B2(new_n516_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT75), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n527_), .A2(new_n533_), .A3(new_n528_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n534_), .A3(new_n523_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536_));
  INV_X1    g335(.A(new_n522_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(KEYINPUT37), .C1(new_n522_), .C2(new_n529_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(G1gat), .ZN(new_n542_));
  INV_X1    g341(.A(G8gat), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT76), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT76), .B(KEYINPUT14), .C1(new_n542_), .C2(new_n543_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G8gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n555_));
  XOR2_X1   g354(.A(G71gat), .B(G78gat), .Z(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n555_), .A2(new_n556_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n553_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G183gat), .B(G211gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n561_), .A2(KEYINPUT17), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(KEYINPUT17), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n561_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n541_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n551_), .A2(new_n461_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n498_), .A2(new_n551_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n551_), .A2(new_n461_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n578_), .B2(new_n572_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G113gat), .B(G141gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT78), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G169gat), .B(G197gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n580_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT71), .ZN(new_n587_));
  XOR2_X1   g386(.A(G120gat), .B(G148gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  INV_X1    g392(.A(new_n560_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n504_), .B2(new_n453_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT69), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n593_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(KEYINPUT69), .B(KEYINPUT12), .C1(new_n495_), .C2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n504_), .A2(new_n453_), .A3(new_n594_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n453_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n560_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n606_), .B2(new_n600_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n592_), .B1(new_n604_), .B2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n602_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n592_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n610_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n587_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n604_), .A2(new_n608_), .A3(new_n592_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n611_), .B1(new_n610_), .B2(new_n607_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(KEYINPUT71), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT13), .ZN(new_n618_));
  AND4_X1   g417(.A1(new_n429_), .A2(new_n571_), .A3(new_n586_), .A4(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n413_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n542_), .A3(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n535_), .A2(new_n537_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n618_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n570_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n586_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n429_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n413_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(new_n385_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n619_), .A2(new_n543_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT103), .B1(new_n629_), .B2(new_n385_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(G8gat), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n629_), .A2(KEYINPUT103), .A3(new_n385_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n636_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AND4_X1   g439(.A1(new_n636_), .A2(new_n639_), .A3(G8gat), .A4(new_n637_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT40), .B(new_n635_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1325gat));
  OAI21_X1  g445(.A(G15gat), .B1(new_n629_), .B2(new_n327_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT41), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n619_), .A2(new_n319_), .A3(new_n386_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1326gat));
  XOR2_X1   g449(.A(new_n281_), .B(KEYINPUT104), .Z(new_n651_));
  OAI21_X1  g450(.A(G22gat), .B1(new_n629_), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT42), .ZN(new_n653_));
  INV_X1    g452(.A(G22gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n651_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n619_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n624_), .A2(new_n570_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n429_), .A2(new_n586_), .A3(new_n618_), .A4(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n620_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n618_), .A2(new_n626_), .A3(new_n586_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT105), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  INV_X1    g463(.A(new_n541_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n429_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n388_), .A2(new_n413_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n667_), .B2(new_n541_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n663_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT44), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n670_), .A2(G29gat), .A3(new_n620_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n664_), .B1(new_n429_), .B2(new_n665_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n667_), .A2(KEYINPUT43), .A3(new_n541_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n675_), .B2(new_n663_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n661_), .B1(new_n671_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n385_), .A2(G36gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT107), .B1(new_n659_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n659_), .A2(KEYINPUT107), .A3(new_n683_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n686_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT45), .B1(new_n689_), .B2(new_n684_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n385_), .B1(new_n669_), .B2(KEYINPUT44), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n679_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n681_), .B1(new_n691_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n677_), .B1(new_n669_), .B2(KEYINPUT106), .ZN(new_n696_));
  AOI211_X1 g495(.A(new_n672_), .B(new_n663_), .C1(new_n666_), .C2(new_n668_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n693_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G36gat), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n688_), .A2(new_n690_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n695_), .A2(new_n702_), .ZN(G1329gat));
  NOR3_X1   g502(.A1(new_n659_), .A2(G43gat), .A3(new_n327_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n327_), .B1(new_n669_), .B2(KEYINPUT44), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n706_), .B2(G43gat), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT47), .B(new_n704_), .C1(new_n706_), .C2(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n660_), .B2(new_n655_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n670_), .A2(G50gat), .A3(new_n281_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n679_), .ZN(G1331gat));
  NOR3_X1   g513(.A1(new_n618_), .A2(new_n626_), .A3(new_n586_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n429_), .A2(new_n624_), .A3(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n413_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n429_), .A2(new_n571_), .A3(new_n627_), .A4(new_n625_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n413_), .A2(G57gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT108), .Z(G1332gat));
  OAI21_X1  g520(.A(G64gat), .B1(new_n716_), .B2(new_n385_), .ZN(new_n722_));
  XOR2_X1   g521(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n385_), .A2(G64gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n718_), .B2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n716_), .B2(new_n327_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n327_), .A2(G71gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n718_), .B2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n716_), .B2(new_n651_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n651_), .A2(G78gat), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT110), .Z(new_n734_));
  OR2_X1    g533(.A1(new_n734_), .A2(new_n718_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT111), .ZN(G1335gat));
  AND4_X1   g536(.A1(new_n429_), .A2(new_n627_), .A3(new_n625_), .A4(new_n658_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n440_), .A3(new_n620_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT112), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n744_), .A2(KEYINPUT113), .A3(new_n746_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n620_), .A3(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n739_), .B1(new_n751_), .B2(new_n440_), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n738_), .B2(new_n634_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n749_), .A2(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n634_), .A2(new_n490_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT114), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n754_), .B2(new_n756_), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n738_), .A2(new_n386_), .A3(new_n433_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n327_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n469_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g560(.A1(new_n738_), .A2(new_n434_), .A3(new_n281_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n745_), .A2(new_n281_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G106gat), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT52), .B(new_n434_), .C1(new_n745_), .C2(new_n281_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g567(.A1(new_n387_), .A2(new_n413_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT12), .B1(new_n606_), .B2(KEYINPUT69), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n596_), .B(new_n593_), .C1(new_n605_), .C2(new_n560_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n600_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT117), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n599_), .A2(new_n775_), .A3(new_n600_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n601_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n778_));
  NOR2_X1   g577(.A1(new_n610_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(KEYINPUT55), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n602_), .B(new_n782_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n779_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT56), .B(new_n611_), .C1(new_n777_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n611_), .B1(new_n777_), .B2(new_n784_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n601_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n775_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n600_), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT117), .B(new_n793_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n610_), .A2(new_n781_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n610_), .B2(new_n778_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n611_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n790_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n580_), .A2(new_n585_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n573_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n575_), .B1(new_n578_), .B2(new_n572_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n584_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n612_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(KEYINPUT58), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n800_), .A2(new_n806_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n665_), .A2(new_n807_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n586_), .A2(new_n812_), .A3(new_n614_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n586_), .B2(new_n614_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n611_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n789_), .B(new_n592_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  INV_X1    g618(.A(new_n805_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT118), .B1(new_n617_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n822_), .B(new_n805_), .C1(new_n613_), .C2(new_n616_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n818_), .B(new_n819_), .C1(new_n821_), .C2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n535_), .A2(new_n819_), .A3(new_n537_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n811_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT121), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n811_), .B(new_n832_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n626_), .A3(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n541_), .A2(new_n570_), .A3(new_n627_), .A4(new_n618_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT54), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n770_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n586_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n818_), .A2(new_n819_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n821_), .A2(new_n823_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n826_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT57), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT58), .B1(new_n800_), .B2(new_n806_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n541_), .A2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n843_), .A2(new_n827_), .B1(new_n845_), .B2(new_n807_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n836_), .B1(new_n570_), .B2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n770_), .A2(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n586_), .B(new_n849_), .C1(new_n837_), .C2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n839_), .B1(new_n852_), .B2(new_n838_), .ZN(G1340gat));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n626_), .B1(new_n846_), .B2(new_n832_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n833_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n836_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n850_), .B1(new_n857_), .B2(new_n769_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n849_), .A2(new_n625_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n854_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n618_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT123), .B(new_n861_), .C1(new_n837_), .C2(new_n850_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(G120gat), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G120gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(G120gat), .B1(new_n625_), .B2(new_n864_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n867_), .B2(new_n866_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n837_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n863_), .A2(new_n870_), .ZN(G1341gat));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n837_), .A2(new_n872_), .A3(new_n570_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n570_), .B(new_n849_), .C1(new_n837_), .C2(new_n850_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(new_n872_), .ZN(G1342gat));
  OAI21_X1  g675(.A(new_n849_), .B1(new_n837_), .B2(new_n850_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G134gat), .B1(new_n877_), .B2(new_n541_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n837_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n624_), .A2(G134gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n281_), .A2(new_n327_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n882_), .A2(new_n413_), .A3(new_n634_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n857_), .A2(new_n586_), .A3(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n857_), .A2(new_n625_), .A3(new_n883_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g686(.A1(new_n857_), .A2(new_n570_), .A3(new_n883_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  NOR2_X1   g689(.A1(new_n624_), .A2(G162gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n857_), .A2(new_n883_), .A3(new_n891_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n857_), .A2(new_n665_), .A3(new_n883_), .ZN(new_n893_));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n847_), .A2(new_n651_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n620_), .A2(new_n327_), .A3(new_n385_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n897_), .A2(new_n334_), .A3(new_n586_), .A4(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n586_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT124), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n903_), .B2(G169gat), .ZN(new_n904_));
  AOI211_X1 g703(.A(KEYINPUT62), .B(new_n311_), .C1(new_n897_), .C2(new_n902_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n899_), .B1(new_n904_), .B2(new_n905_), .ZN(G1348gat));
  INV_X1    g705(.A(new_n898_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n896_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G176gat), .B1(new_n908_), .B2(new_n625_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n281_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n907_), .A2(new_n312_), .A3(new_n618_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(G1349gat));
  NOR2_X1   g711(.A1(new_n907_), .A2(new_n626_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n896_), .A2(new_n308_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n910_), .A2(new_n913_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n916_), .B(KEYINPUT125), .C1(new_n917_), .C2(G183gat), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n910_), .B2(new_n913_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n915_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n921_), .ZN(G1350gat));
  NAND4_X1  g721(.A1(new_n908_), .A2(new_n309_), .A3(new_n537_), .A4(new_n535_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n896_), .A2(new_n541_), .A3(new_n907_), .ZN(new_n924_));
  INV_X1    g723(.A(G190gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n620_), .A2(new_n882_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT126), .Z(new_n928_));
  NAND3_X1  g727(.A1(new_n857_), .A2(new_n634_), .A3(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n627_), .ZN(new_n930_));
  INV_X1    g729(.A(G197gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n929_), .A2(new_n618_), .ZN(new_n933_));
  INV_X1    g732(.A(G204gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1353gat));
  AOI21_X1  g734(.A(new_n626_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n929_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT127), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n938_), .B(new_n941_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n929_), .B2(new_n541_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n624_), .A2(G218gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n929_), .B2(new_n944_), .ZN(G1355gat));
endmodule


