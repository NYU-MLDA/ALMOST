//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n204_), .B(new_n205_), .C1(G183gat), .C2(G190gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n207_));
  OR3_X1    g006(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n204_), .A2(new_n205_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n214_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n216_), .B(new_n217_), .C1(new_n219_), .C2(KEYINPUT24), .ZN(new_n220_));
  INV_X1    g019(.A(G190gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT26), .B1(new_n221_), .B2(KEYINPUT77), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(G183gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT25), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n222_), .B(new_n225_), .C1(KEYINPUT76), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(KEYINPUT76), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n226_), .A2(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n209_), .B1(new_n220_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G197gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G204gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT21), .B1(new_n235_), .B2(KEYINPUT88), .ZN(new_n236_));
  INV_X1    g035(.A(G204gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G197gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n236_), .B1(new_n240_), .B2(KEYINPUT88), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n239_), .B2(KEYINPUT21), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(KEYINPUT21), .ZN(new_n244_));
  OAI22_X1  g043(.A1(new_n241_), .A2(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n233_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT95), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT19), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT20), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(G169gat), .B2(G176gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n219_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n218_), .A2(new_n253_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n230_), .A3(new_n227_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n255_), .A2(new_n217_), .A3(new_n256_), .A4(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT22), .B(G169gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n212_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n215_), .B(KEYINPUT92), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n206_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT93), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n264_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n259_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n248_), .B(new_n252_), .C1(new_n245_), .C2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT20), .B1(new_n233_), .B2(new_n245_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT90), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n245_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT90), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n272_), .B(KEYINPUT20), .C1(new_n233_), .C2(new_n245_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(KEYINPUT94), .A3(new_n250_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT94), .B1(new_n274_), .B2(new_n250_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n268_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G8gat), .B(G36gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT97), .ZN(new_n285_));
  INV_X1    g084(.A(new_n283_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n286_), .B(new_n268_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n276_), .A2(new_n277_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n290_), .A2(KEYINPUT97), .A3(new_n286_), .A4(new_n268_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n287_), .A2(KEYINPUT100), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(KEYINPUT100), .ZN(new_n294_));
  INV_X1    g093(.A(new_n274_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n263_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n245_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n251_), .B1(new_n297_), .B2(new_n259_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n248_), .A2(new_n298_), .ZN(new_n299_));
  MUX2_X1   g098(.A(new_n295_), .B(new_n299_), .S(new_n250_), .Z(new_n300_));
  AOI21_X1  g099(.A(new_n289_), .B1(new_n300_), .B2(new_n283_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n293_), .A2(new_n294_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n292_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT1), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT86), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309_));
  INV_X1    g108(.A(G155gat), .ZN(new_n310_));
  INV_X1    g109(.A(G162gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(KEYINPUT1), .B2(new_n306_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n304_), .B(new_n305_), .C1(new_n308_), .C2(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n305_), .A2(KEYINPUT3), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n304_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n305_), .A2(KEYINPUT3), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .A4(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(new_n306_), .A3(new_n314_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT29), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n325_), .B(KEYINPUT28), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(KEYINPUT29), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n245_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n326_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT89), .ZN(new_n331_));
  INV_X1    g130(.A(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(G228gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(G228gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n331_), .B(new_n336_), .Z(new_n337_));
  XOR2_X1   g136(.A(G22gat), .B(G50gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n328_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n326_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n339_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350_));
  OR3_X1    g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n324_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n316_), .A2(new_n351_), .A3(new_n323_), .A4(new_n352_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT4), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n358_), .C1(KEYINPUT4), .C2(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n355_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT98), .B1(new_n360_), .B2(new_n358_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT98), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n354_), .A2(new_n362_), .A3(new_n357_), .A4(new_n355_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G85gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n359_), .A2(new_n368_), .A3(new_n361_), .A4(new_n363_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n233_), .B(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n374_), .A2(KEYINPUT82), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(KEYINPUT82), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G71gat), .B(G99gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT80), .B(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT81), .B(G15gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n380_), .B(new_n383_), .Z(new_n384_));
  NOR2_X1   g183(.A1(new_n377_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n375_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n353_), .B(KEYINPUT84), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(KEYINPUT31), .Z(new_n389_));
  OR3_X1    g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n389_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n372_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n303_), .A2(KEYINPUT101), .A3(new_n345_), .A4(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n292_), .A2(new_n302_), .A3(new_n345_), .A4(new_n392_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT101), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n345_), .A2(new_n372_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n292_), .A2(new_n397_), .A3(new_n302_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n286_), .A2(KEYINPUT32), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n300_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n372_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n278_), .A2(new_n399_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n288_), .A2(new_n291_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT99), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n371_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n371_), .B2(new_n406_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n356_), .B1(KEYINPUT4), .B2(new_n354_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(new_n358_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n369_), .B1(new_n360_), .B2(new_n357_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT33), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n407_), .A2(new_n408_), .B1(new_n371_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n403_), .B1(new_n404_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n345_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n398_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n390_), .A2(new_n391_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n393_), .A2(new_n396_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G120gat), .B(G148gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT5), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G176gat), .B(G204gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  XOR2_X1   g222(.A(new_n423_), .B(KEYINPUT68), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT66), .ZN(new_n426_));
  INV_X1    g225(.A(G85gat), .ZN(new_n427_));
  INV_X1    g226(.A(G92gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT65), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G92gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n426_), .B1(new_n432_), .B2(KEYINPUT9), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT9), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT65), .B(G92gat), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT66), .B(new_n434_), .C1(new_n435_), .C2(new_n427_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n427_), .A2(new_n428_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n438_), .B2(KEYINPUT9), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n433_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT67), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT67), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n433_), .A2(new_n442_), .A3(new_n436_), .A4(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT10), .B(G99gat), .ZN(new_n447_));
  OR3_X1    g246(.A1(new_n447_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT64), .B1(new_n447_), .B2(G106gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n446_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n441_), .A2(new_n443_), .A3(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n438_), .A2(new_n437_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT7), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n452_), .B1(new_n455_), .B2(new_n446_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT8), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n460_));
  XOR2_X1   g259(.A(G71gat), .B(G78gat), .Z(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n461_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n458_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n451_), .A2(new_n457_), .A3(new_n466_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT12), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n466_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G230gat), .A2(G233gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n425_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(new_n477_), .B(new_n423_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT13), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT13), .B1(new_n479_), .B2(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G229gat), .A2(G233gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G15gat), .B(G22gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(G1gat), .A2(G8gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(KEYINPUT14), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT72), .ZN(new_n491_));
  XOR2_X1   g290(.A(G1gat), .B(G8gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n490_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n499_), .A2(KEYINPUT69), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(KEYINPUT69), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n501_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n502_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n498_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n493_), .A2(new_n497_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n503_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n487_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n509_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n506_), .A2(KEYINPUT15), .A3(new_n503_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n498_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n512_), .A2(new_n517_), .A3(new_n486_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  NAND3_X1  g320(.A1(new_n511_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n511_), .B2(new_n518_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n485_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n419_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT34), .Z(new_n529_));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n458_), .A2(new_n515_), .A3(new_n514_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n531_), .B1(new_n532_), .B2(KEYINPUT70), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n516_), .A2(new_n458_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n451_), .A2(new_n509_), .A3(new_n457_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n530_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n534_), .A2(KEYINPUT70), .A3(new_n531_), .A4(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G190gat), .B(G218gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT71), .B1(new_n538_), .B2(new_n539_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT36), .B1(new_n549_), .B2(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n540_), .A2(new_n546_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT37), .A4(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT73), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n466_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n498_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G127gat), .B(G155gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n561_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT75), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n566_), .A2(new_n567_), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n561_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n557_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n527_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT102), .Z(new_n576_));
  INV_X1    g375(.A(G1gat), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n372_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT38), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n393_), .A2(new_n396_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n416_), .A2(new_n418_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n552_), .B(KEYINPUT103), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n526_), .A2(new_n573_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT104), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(KEYINPUT104), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n372_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT105), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT105), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n580_), .B(new_n581_), .C1(new_n594_), .C2(new_n595_), .ZN(G1324gat));
  INV_X1    g395(.A(G8gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n303_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n576_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G8gat), .B1(new_n587_), .B2(new_n303_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT106), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(KEYINPUT106), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n599_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(KEYINPUT40), .B(new_n599_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1325gat));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n576_), .A2(new_n611_), .A3(new_n417_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n590_), .A2(new_n417_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n613_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(new_n613_), .B2(G15gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(G1326gat));
  NOR2_X1   g415(.A1(new_n345_), .A2(G22gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT108), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n576_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(G22gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n590_), .B2(new_n415_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n619_), .B1(new_n623_), .B2(new_n624_), .ZN(G1327gat));
  INV_X1    g424(.A(new_n552_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n573_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n527_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(G29gat), .B1(new_n629_), .B2(new_n372_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n419_), .B2(new_n556_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n394_), .B(KEYINPUT101), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n407_), .A2(new_n408_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n412_), .A2(new_n371_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n291_), .B2(new_n288_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n345_), .B1(new_n637_), .B2(new_n403_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n417_), .B1(new_n638_), .B2(new_n398_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n632_), .B(new_n557_), .C1(new_n633_), .C2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n631_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n526_), .A2(new_n627_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(KEYINPUT44), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT44), .B1(new_n641_), .B2(new_n642_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n372_), .A2(G29gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n630_), .B1(new_n645_), .B2(new_n646_), .ZN(G1328gat));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n643_), .A2(new_n644_), .A3(new_n303_), .ZN(new_n649_));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n629_), .A2(new_n650_), .A3(new_n598_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT45), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n652_), .B(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(KEYINPUT46), .C1(new_n650_), .C2(new_n649_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(G1329gat));
  AOI21_X1  g457(.A(G43gat), .B1(new_n629_), .B2(new_n417_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT109), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n645_), .A2(G43gat), .A3(new_n417_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1330gat));
  AOI21_X1  g466(.A(G50gat), .B1(new_n629_), .B2(new_n415_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n415_), .A2(G50gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n645_), .B2(new_n669_), .ZN(G1331gat));
  INV_X1    g469(.A(new_n485_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n523_), .A2(new_n524_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n584_), .A2(new_n585_), .A3(new_n671_), .A4(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G57gat), .B1(new_n675_), .B2(new_n592_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT111), .B1(new_n584_), .B2(new_n672_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n485_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n584_), .A2(KEYINPUT111), .A3(new_n672_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n574_), .A3(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n592_), .A2(G57gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n676_), .B1(new_n680_), .B2(new_n681_), .ZN(G1332gat));
  OAI21_X1  g481(.A(G64gat), .B1(new_n675_), .B2(new_n303_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT48), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n303_), .A2(G64gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n680_), .B2(new_n685_), .ZN(G1333gat));
  OAI21_X1  g485(.A(G71gat), .B1(new_n675_), .B2(new_n418_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT49), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n418_), .A2(G71gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n680_), .B2(new_n689_), .ZN(G1334gat));
  OAI21_X1  g489(.A(G78gat), .B1(new_n675_), .B2(new_n345_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT50), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n345_), .A2(G78gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n680_), .B2(new_n693_), .ZN(G1335gat));
  NAND3_X1  g493(.A1(new_n678_), .A2(new_n628_), .A3(new_n679_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n372_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n485_), .A2(new_n627_), .A3(new_n525_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n641_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT112), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n592_), .A2(new_n427_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1336gat));
  AOI21_X1  g501(.A(G92gat), .B1(new_n696_), .B2(new_n598_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n303_), .A2(new_n435_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n700_), .B2(new_n704_), .ZN(G1337gat));
  NOR2_X1   g504(.A1(new_n418_), .A2(new_n447_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n698_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n631_), .B2(new_n640_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n417_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n696_), .A2(new_n706_), .B1(G99gat), .B2(new_n709_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g510(.A(G106gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n696_), .A2(new_n712_), .A3(new_n415_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n345_), .B(new_n707_), .C1(new_n631_), .C2(new_n640_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n708_), .B2(new_n415_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n714_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n641_), .A2(new_n716_), .A3(new_n415_), .A4(new_n698_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G106gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(KEYINPUT52), .A3(new_n718_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n713_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT53), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(new_n713_), .C1(new_n720_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1339gat));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT54), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n674_), .A2(new_n485_), .A3(KEYINPUT114), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n556_), .A4(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT115), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n556_), .A2(new_n732_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n673_), .B1(new_n484_), .B2(new_n483_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(KEYINPUT114), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT54), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n736_), .A2(KEYINPUT114), .B1(new_n554_), .B2(new_n555_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT115), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n731_), .A4(new_n730_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n734_), .A2(new_n738_), .A3(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n743_));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n672_), .A2(new_n480_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n475_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n470_), .A2(new_n746_), .A3(new_n473_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n476_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n474_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n475_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n451_), .A2(new_n457_), .A3(new_n466_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n751_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n473_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT55), .B(new_n475_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n749_), .A2(new_n750_), .A3(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n424_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n424_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n745_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n486_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n521_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n512_), .A2(new_n517_), .A3(new_n487_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n522_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n481_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n744_), .B1(new_n768_), .B2(new_n626_), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT117), .B(new_n552_), .C1(new_n760_), .C2(new_n767_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n743_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n765_), .A2(new_n480_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT58), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT58), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n772_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n557_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n556_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT119), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n552_), .B1(new_n760_), .B2(new_n767_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT57), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n771_), .A2(new_n780_), .A3(new_n782_), .A4(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n742_), .B1(new_n785_), .B2(new_n573_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n598_), .A2(new_n415_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n418_), .A2(new_n592_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT59), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(G113gat), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n672_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT121), .ZN(new_n793_));
  INV_X1    g592(.A(new_n743_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n480_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n525_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n757_), .A2(new_n424_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n424_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n626_), .B1(new_n801_), .B2(new_n766_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT117), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n783_), .A2(new_n744_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n794_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n793_), .B1(new_n805_), .B2(new_n781_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n771_), .A2(KEYINPUT121), .A3(new_n778_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n784_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n742_), .B1(new_n808_), .B2(new_n573_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n789_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n810_), .A2(KEYINPUT120), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(KEYINPUT120), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n790_), .B(new_n792_), .C1(new_n809_), .C2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n784_), .B1(new_n781_), .B2(KEYINPUT119), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n779_), .B(new_n556_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n627_), .B1(new_n818_), .B2(new_n771_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n810_), .B1(new_n819_), .B2(new_n742_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n791_), .B1(new_n820_), .B2(new_n672_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n815_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n815_), .A2(KEYINPUT122), .A3(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n485_), .B1(new_n820_), .B2(KEYINPUT59), .ZN(new_n828_));
  INV_X1    g627(.A(new_n814_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n784_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n771_), .A2(new_n778_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n793_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n627_), .B1(new_n832_), .B2(new_n807_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n833_), .B2(new_n742_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n827_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n820_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n827_), .B1(new_n485_), .B2(KEYINPUT60), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n827_), .A2(KEYINPUT60), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT123), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n790_), .A2(new_n671_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n808_), .A2(new_n573_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n742_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n814_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G120gat), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n840_), .A2(new_n848_), .ZN(G1341gat));
  NAND2_X1  g648(.A1(new_n834_), .A2(new_n790_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G127gat), .B1(new_n850_), .B2(new_n573_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n573_), .A2(G127gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n820_), .B2(new_n852_), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n850_), .B2(new_n556_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n585_), .A2(G134gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n820_), .B2(new_n855_), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n786_), .A2(new_n417_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n598_), .A2(new_n592_), .A3(new_n345_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n672_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT124), .B(G141gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n671_), .A3(new_n858_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g663(.A1(new_n859_), .A2(new_n573_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  OAI21_X1  g666(.A(G162gat), .B1(new_n859_), .B2(new_n556_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n585_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n311_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n859_), .B2(new_n870_), .ZN(G1347gat));
  NAND2_X1  g670(.A1(new_n598_), .A2(new_n392_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT125), .Z(new_n873_));
  OR2_X1    g672(.A1(new_n873_), .A2(new_n415_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n809_), .A2(new_n672_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n211_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(new_n211_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n260_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(G1348gat));
  NOR2_X1   g679(.A1(new_n809_), .A2(new_n874_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G176gat), .B1(new_n881_), .B2(new_n671_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n786_), .A2(new_n415_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n873_), .A2(new_n212_), .A3(new_n485_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1349gat));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n230_), .A2(new_n227_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n627_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n886_), .B1(new_n881_), .B2(new_n889_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n809_), .A2(KEYINPUT126), .A3(new_n874_), .A4(new_n888_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n873_), .A2(new_n573_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G183gat), .B1(new_n883_), .B2(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n890_), .A2(new_n891_), .A3(new_n893_), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n881_), .A2(new_n869_), .A3(new_n257_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n809_), .A2(new_n556_), .A3(new_n874_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n221_), .ZN(G1351gat));
  NOR3_X1   g696(.A1(new_n303_), .A2(new_n372_), .A3(new_n345_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n857_), .A2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n672_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n234_), .ZN(G1352gat));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n485_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(new_n237_), .ZN(G1353gat));
  XNOR2_X1  g702(.A(KEYINPUT63), .B(G211gat), .ZN(new_n904_));
  OR2_X1    g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n857_), .A2(new_n627_), .A3(new_n898_), .ZN(new_n906_));
  MUX2_X1   g705(.A(new_n904_), .B(new_n905_), .S(new_n906_), .Z(G1354gat));
  INV_X1    g706(.A(G218gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n899_), .A2(new_n908_), .A3(new_n556_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n899_), .A2(new_n585_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  AOI21_X1  g710(.A(G218gat), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT127), .B1(new_n899_), .B2(new_n585_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n909_), .B1(new_n912_), .B2(new_n913_), .ZN(G1355gat));
endmodule


