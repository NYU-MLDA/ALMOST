//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n971_, new_n972_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n984_;
  XNOR2_X1  g000(.A(G1gat), .B(G8gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G15gat), .ZN(new_n205_));
  INV_X1    g004(.A(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G15gat), .A2(G22gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G1gat), .A2(G8gat), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n207_), .A2(new_n208_), .B1(KEYINPUT14), .B2(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n204_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n204_), .A2(new_n210_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT75), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n214_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n217_), .A2(new_n221_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n204_), .B(new_n210_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n222_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n213_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n230_), .A3(new_n226_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G169gat), .B(G197gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  AND3_X1   g038(.A1(new_n232_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G8gat), .B(G36gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT18), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G64gat), .B(G92gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT19), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT93), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT85), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT82), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT82), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(G169gat), .A3(G176gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G183gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT25), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G183gat), .ZN(new_n263_));
  INV_X1    g062(.A(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT26), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT26), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G190gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n261_), .A2(new_n263_), .A3(new_n265_), .A4(new_n267_), .ZN(new_n268_));
  OR3_X1    g067(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n259_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT23), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n273_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n270_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G169gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT22), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT22), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G169gat), .ZN(new_n284_));
  INV_X1    g083(.A(G176gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n275_), .A2(KEYINPUT23), .A3(new_n276_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n278_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n271_), .B2(KEYINPUT23), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n287_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n252_), .B1(new_n280_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n276_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT83), .B1(G183gat), .B2(G190gat), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n278_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n291_), .A2(new_n289_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n294_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n287_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n278_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n272_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n305_), .A2(new_n259_), .A3(new_n269_), .A4(new_n268_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n306_), .A3(KEYINPUT85), .ZN(new_n307_));
  XOR2_X1   g106(.A(G197gat), .B(G204gat), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n310_), .A2(new_n313_), .A3(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n296_), .A2(new_n307_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n251_), .B1(new_n318_), .B2(KEYINPUT20), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n282_), .A2(new_n284_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(KEYINPUT97), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n285_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n256_), .A2(new_n258_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n305_), .A2(new_n294_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n266_), .A2(G190gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n264_), .A2(KEYINPUT26), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n261_), .A2(new_n263_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n265_), .A2(new_n267_), .A3(KEYINPUT94), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n254_), .A2(new_n255_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(KEYINPUT95), .A3(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n292_), .A2(new_n269_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT96), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n333_), .A2(KEYINPUT95), .A3(new_n334_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT95), .B1(new_n333_), .B2(new_n334_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT96), .B(new_n341_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n326_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n319_), .B1(new_n347_), .B2(new_n316_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n318_), .A2(new_n251_), .A3(KEYINPUT20), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n250_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n326_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT96), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n354_), .B2(new_n345_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n317_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n317_), .B1(new_n296_), .B2(new_n307_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n249_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n247_), .B1(new_n350_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n318_), .A2(KEYINPUT20), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT93), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(new_n349_), .C1(new_n317_), .C2(new_n355_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n249_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n246_), .A3(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n365_), .A2(new_n249_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n246_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n246_), .B(KEYINPUT103), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n365_), .A2(new_n249_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n326_), .A2(new_n352_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n316_), .B1(new_n374_), .B2(KEYINPUT100), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(KEYINPUT100), .B2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n357_), .A2(new_n358_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n250_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n372_), .B1(new_n373_), .B2(new_n378_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n368_), .A2(new_n369_), .B1(new_n371_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  AND2_X1   g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT1), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  OAI22_X1  g185(.A1(new_n385_), .A2(KEYINPUT89), .B1(new_n386_), .B2(KEYINPUT1), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT89), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n388_), .A3(new_n383_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n384_), .A2(new_n387_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G141gat), .B(G148gat), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n394_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(KEYINPUT3), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n394_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n382_), .A2(new_n385_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n393_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G134gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G127gat), .ZN(new_n407_));
  INV_X1    g206(.A(G127gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G134gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G120gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G113gat), .ZN(new_n412_));
  INV_X1    g211(.A(G113gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G120gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .A4(new_n414_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT87), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n410_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n412_), .A4(new_n414_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n405_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(new_n417_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n393_), .A2(new_n404_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT99), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n423_), .A2(KEYINPUT4), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n418_), .A2(new_n421_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n391_), .A2(new_n392_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n425_), .B(KEYINPUT4), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT98), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n423_), .A2(KEYINPUT98), .A3(KEYINPUT4), .A4(new_n425_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n430_), .B1(new_n438_), .B2(new_n429_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G85gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT0), .B(G57gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(new_n430_), .C1(new_n438_), .C2(new_n429_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(KEYINPUT101), .A3(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n438_), .A2(new_n429_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n445_), .A4(new_n430_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT102), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n447_), .A2(new_n450_), .A3(KEYINPUT102), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n296_), .A2(new_n307_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT86), .B(G43gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n456_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(new_n422_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(new_n205_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT30), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT31), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n461_), .B(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT28), .ZN(new_n468_));
  XOR2_X1   g267(.A(G22gat), .B(G50gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n471_));
  OAI21_X1  g270(.A(G78gat), .B1(new_n471_), .B2(new_n317_), .ZN(new_n472_));
  INV_X1    g271(.A(G78gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n473_), .B(new_n316_), .C1(new_n433_), .C2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(G106gat), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(G106gat), .A3(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G228gat), .A2(G233gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT91), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n317_), .B2(KEYINPUT92), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n478_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n481_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n478_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n476_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n470_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n470_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n380_), .A2(new_n455_), .A3(new_n466_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n482_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n470_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n486_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n380_), .A2(new_n455_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n444_), .A2(KEYINPUT33), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT33), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n439_), .A2(new_n498_), .A3(new_n443_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n438_), .A2(new_n429_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n501_), .B(new_n445_), .C1(new_n429_), .C2(new_n426_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n500_), .A2(new_n362_), .A3(new_n367_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n246_), .A2(KEYINPUT32), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n373_), .B2(new_n378_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n366_), .A2(new_n360_), .A3(new_n504_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(new_n450_), .A3(new_n447_), .A4(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n489_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n466_), .B1(new_n496_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT104), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n491_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n489_), .B1(new_n454_), .B2(new_n453_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n514_), .A2(new_n380_), .B1(new_n509_), .B2(new_n489_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT104), .B1(new_n515_), .B2(new_n466_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n242_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT67), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT66), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT11), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G71gat), .B(G78gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n518_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  AOI211_X1 g324(.A(KEYINPUT67), .B(new_n523_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n526_));
  OAI22_X1  g325(.A1(new_n525_), .A2(new_n526_), .B1(new_n521_), .B2(new_n520_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT66), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n519_), .B(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT67), .B1(new_n530_), .B2(new_n523_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n522_), .A2(new_n518_), .A3(new_n524_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n520_), .A2(new_n521_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G99gat), .ZN(new_n535_));
  INV_X1    g334(.A(G106gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT6), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT6), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT64), .ZN(new_n541_));
  XOR2_X1   g340(.A(G85gat), .B(G92gat), .Z(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT9), .ZN(new_n543_));
  INV_X1    g342(.A(G85gat), .ZN(new_n544_));
  INV_X1    g343(.A(G92gat), .ZN(new_n545_));
  OR3_X1    g344(.A1(new_n544_), .A2(new_n545_), .A3(KEYINPUT9), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT10), .B(G99gat), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n543_), .B(new_n546_), .C1(G106gat), .C2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n541_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT8), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT65), .ZN(new_n552_));
  NOR2_X1   g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n550_), .B(new_n542_), .C1(new_n541_), .C2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n540_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n550_), .B1(new_n557_), .B2(new_n542_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n549_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n527_), .A2(new_n534_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n527_), .B2(new_n534_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n527_), .A2(new_n534_), .A3(new_n560_), .A4(KEYINPUT68), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n563_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G230gat), .A2(G233gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n561_), .A2(new_n568_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT12), .B1(new_n560_), .B2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n564_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n564_), .A2(new_n573_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G120gat), .B(G148gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT71), .ZN(new_n578_));
  XOR2_X1   g377(.A(G176gat), .B(G204gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n570_), .A2(new_n576_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT72), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n564_), .B(new_n573_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n585_), .A2(new_n571_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n582_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n586_), .A2(new_n582_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(KEYINPUT13), .A3(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(G231gat), .ZN(new_n597_));
  INV_X1    g396(.A(G233gat), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n527_), .A2(new_n534_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n600_), .A2(KEYINPUT80), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(KEYINPUT80), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n599_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n601_), .A2(new_n602_), .A3(new_n599_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n604_), .A2(new_n225_), .A3(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n225_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT16), .ZN(new_n610_));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n572_), .A3(KEYINPUT17), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n614_), .B1(KEYINPUT17), .B2(new_n613_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n606_), .A2(new_n607_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n222_), .B(KEYINPUT15), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n560_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n560_), .A2(new_n224_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n542_), .A2(new_n550_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT64), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n540_), .B(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n633_), .B2(new_n554_), .ZN(new_n634_));
  OAI22_X1  g433(.A1(new_n634_), .A2(new_n558_), .B1(new_n541_), .B2(new_n548_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n234_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n624_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n628_), .A4(new_n627_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n630_), .A2(KEYINPUT78), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640_));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641_));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n640_), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n630_), .A2(new_n645_), .A3(new_n638_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n640_), .B1(new_n639_), .B2(new_n646_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n618_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n639_), .A2(new_n646_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT36), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n653_), .A2(KEYINPUT37), .A3(new_n648_), .A4(new_n647_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n615_), .A2(new_n617_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n517_), .A2(new_n596_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT105), .ZN(new_n657_));
  INV_X1    g456(.A(G1gat), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n447_), .A2(KEYINPUT102), .A3(new_n450_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT102), .B1(new_n447_), .B2(new_n450_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n657_), .A2(KEYINPUT38), .A3(new_n658_), .A4(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n232_), .A2(new_n236_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n239_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n232_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n671_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n653_), .A2(KEYINPUT106), .A3(new_n648_), .A4(new_n647_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n615_), .A2(new_n617_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AND4_X1   g476(.A1(new_n670_), .A2(new_n675_), .A3(new_n596_), .A4(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n661_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G1gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n664_), .A2(new_n665_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n664_), .A2(KEYINPUT107), .A3(new_n665_), .A4(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1324gat));
  INV_X1    g484(.A(G8gat), .ZN(new_n686_));
  AOI221_X4 g485(.A(new_n247_), .B1(new_n356_), .B2(new_n359_), .C1(new_n365_), .C2(new_n249_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n246_), .B1(new_n366_), .B2(new_n360_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n369_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n379_), .A2(KEYINPUT27), .A3(new_n367_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n657_), .A2(new_n686_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n678_), .A2(new_n691_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(G8gat), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n693_), .B2(G8gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g497(.A1(new_n657_), .A2(new_n205_), .A3(new_n466_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n678_), .A2(new_n466_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n700_), .B2(G15gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(G1326gat));
  AOI21_X1  g503(.A(new_n206_), .B1(new_n678_), .B2(new_n495_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT42), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n657_), .A2(new_n206_), .A3(new_n495_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1327gat));
  NAND2_X1  g507(.A1(new_n676_), .A2(new_n674_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n517_), .A2(new_n596_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(G29gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n661_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n651_), .A2(new_n654_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n466_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n495_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n691_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n495_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n512_), .B(new_n716_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n490_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n496_), .A2(new_n510_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n512_), .B1(new_n722_), .B2(new_n716_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n715_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT43), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n516_), .A2(new_n490_), .A3(new_n720_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n715_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n677_), .A2(new_n595_), .A3(new_n242_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  INV_X1    g531(.A(new_n730_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n732_), .B(new_n733_), .C1(new_n725_), .C2(new_n728_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n731_), .A2(new_n734_), .A3(new_n455_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n713_), .B1(new_n735_), .B2(new_n712_), .ZN(G1328gat));
  NAND2_X1  g535(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n737_));
  NOR2_X1   g536(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n738_));
  INV_X1    g537(.A(G36gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n711_), .A2(new_n739_), .A3(new_n691_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT45), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n711_), .A2(new_n742_), .A3(new_n739_), .A4(new_n691_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n738_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n731_), .A2(new_n734_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n691_), .ZN(new_n747_));
  AOI211_X1 g546(.A(KEYINPUT43), .B(new_n714_), .C1(new_n513_), .C2(new_n516_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n727_), .B1(new_n726_), .B2(new_n715_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n730_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n732_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT44), .B(new_n730_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n751_), .A2(new_n745_), .A3(new_n691_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G36gat), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n737_), .B(new_n744_), .C1(new_n747_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(new_n691_), .A3(new_n752_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT110), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(G36gat), .A3(new_n753_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n737_), .B1(new_n759_), .B2(new_n744_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n756_), .A2(new_n760_), .ZN(G1329gat));
  NAND2_X1  g560(.A1(new_n746_), .A2(new_n466_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G43gat), .ZN(new_n763_));
  INV_X1    g562(.A(G43gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n711_), .A2(new_n764_), .A3(new_n466_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n763_), .A2(KEYINPUT47), .A3(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1330gat));
  NAND2_X1  g569(.A1(new_n746_), .A2(new_n495_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G50gat), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n489_), .A2(G50gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT112), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n711_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(G1331gat));
  NOR2_X1   g575(.A1(new_n596_), .A2(new_n670_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n726_), .A2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(new_n655_), .ZN(new_n779_));
  INV_X1    g578(.A(G57gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n661_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n675_), .A2(new_n677_), .A3(new_n777_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n783_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(new_n661_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n781_), .B1(new_n787_), .B2(new_n780_), .ZN(G1332gat));
  INV_X1    g587(.A(G64gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(new_n789_), .A3(new_n691_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n691_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G64gat), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(KEYINPUT48), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(KEYINPUT48), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(G1333gat));
  INV_X1    g594(.A(G71gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n796_), .A3(new_n466_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n784_), .A2(new_n466_), .A3(new_n785_), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(G71gat), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G71gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT115), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n797_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1334gat));
  NAND3_X1  g605(.A1(new_n779_), .A2(new_n473_), .A3(new_n495_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n786_), .A2(new_n495_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(G78gat), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(KEYINPUT50), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(KEYINPUT50), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(G1335gat));
  NOR2_X1   g611(.A1(new_n748_), .A2(new_n749_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n729_), .A2(KEYINPUT116), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n596_), .A2(new_n677_), .A3(new_n670_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G85gat), .B1(new_n818_), .B2(new_n455_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n778_), .A2(new_n710_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n544_), .A3(new_n661_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1336gat));
  OAI21_X1  g621(.A(G92gat), .B1(new_n818_), .B2(new_n380_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n545_), .A3(new_n691_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1337gat));
  OAI21_X1  g624(.A(G99gat), .B1(new_n818_), .B2(new_n716_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n547_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n820_), .A2(new_n466_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g629(.A1(new_n817_), .A2(new_n495_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G106gat), .B1(new_n813_), .B2(new_n831_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(KEYINPUT117), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(KEYINPUT117), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(KEYINPUT52), .A3(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n834_), .A2(KEYINPUT52), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n820_), .A2(new_n536_), .A3(new_n495_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT53), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n835_), .A2(new_n836_), .A3(new_n840_), .A4(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1339gat));
  NOR3_X1   g641(.A1(new_n691_), .A2(new_n716_), .A3(new_n495_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n672_), .A2(new_n673_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n587_), .B1(new_n586_), .B2(new_n582_), .ZN(new_n845_));
  AND4_X1   g644(.A1(new_n587_), .A2(new_n570_), .A3(new_n576_), .A4(new_n582_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n670_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT12), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n635_), .B2(KEYINPUT69), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n564_), .B(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n563_), .A2(new_n566_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n569_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n576_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n585_), .A2(KEYINPUT55), .A3(new_n571_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n582_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(KEYINPUT56), .A3(new_n857_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n847_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n239_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n235_), .A2(new_n226_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n231_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n864_), .A2(new_n865_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n863_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n669_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT57), .B(new_n844_), .C1(new_n862_), .C2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT120), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n242_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n856_), .A2(KEYINPUT56), .A3(new_n857_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n857_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n870_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n591_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n674_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n881_), .A3(KEYINPUT57), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n844_), .B1(new_n862_), .B2(new_n871_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n870_), .B1(new_n588_), .B2(new_n584_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n714_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT58), .B(new_n886_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n884_), .A2(new_n885_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n677_), .B1(new_n883_), .B2(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n655_), .A2(new_n242_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n894_));
  OR2_X1    g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(KEYINPUT118), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n661_), .B(new_n843_), .C1(new_n892_), .C2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n413_), .A3(new_n670_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n872_), .A2(KEYINPUT120), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n881_), .B1(new_n880_), .B2(KEYINPUT57), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n891_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n676_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n898_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n455_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n907_), .A2(KEYINPUT121), .A3(KEYINPUT59), .A4(new_n843_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n899_), .B2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n908_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n908_), .B2(new_n911_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n913_), .A2(new_n914_), .A3(new_n242_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n901_), .B1(new_n915_), .B2(new_n413_), .ZN(G1340gat));
  OAI21_X1  g715(.A(new_n411_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n900_), .B(new_n917_), .C1(KEYINPUT60), .C2(new_n411_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n596_), .B1(new_n908_), .B2(new_n911_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n411_), .ZN(G1341gat));
  NAND3_X1  g719(.A1(new_n900_), .A2(new_n408_), .A3(new_n677_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n913_), .A2(new_n914_), .A3(new_n676_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n408_), .ZN(G1342gat));
  NAND3_X1  g722(.A1(new_n900_), .A2(new_n406_), .A3(new_n674_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n913_), .A2(new_n914_), .A3(new_n714_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n406_), .ZN(G1343gat));
  NOR3_X1   g725(.A1(new_n691_), .A2(new_n466_), .A3(new_n489_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n907_), .A2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n670_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n595_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g732(.A1(new_n928_), .A2(new_n676_), .ZN(new_n934_));
  XOR2_X1   g733(.A(KEYINPUT61), .B(G155gat), .Z(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1346gat));
  INV_X1    g735(.A(G162gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n929_), .A2(new_n937_), .A3(new_n674_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n928_), .A2(new_n714_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(KEYINPUT123), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n938_), .B(new_n942_), .C1(new_n937_), .C2(new_n939_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1347gat));
  NAND2_X1  g743(.A1(new_n905_), .A2(new_n906_), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n380_), .A2(new_n661_), .A3(new_n716_), .A4(new_n495_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  OR3_X1    g746(.A1(new_n947_), .A2(KEYINPUT124), .A3(new_n242_), .ZN(new_n948_));
  OAI21_X1  g747(.A(KEYINPUT124), .B1(new_n947_), .B2(new_n242_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n948_), .A2(G169gat), .A3(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n947_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n953_), .A2(new_n321_), .A3(new_n670_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n948_), .A2(KEYINPUT62), .A3(new_n949_), .A4(G169gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n952_), .A2(new_n954_), .A3(new_n955_), .ZN(G1348gat));
  XNOR2_X1  g755(.A(KEYINPUT125), .B(G176gat), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n285_), .A2(KEYINPUT125), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n953_), .A2(new_n595_), .ZN(new_n959_));
  MUX2_X1   g758(.A(new_n957_), .B(new_n958_), .S(new_n959_), .Z(G1349gat));
  OAI21_X1  g759(.A(new_n260_), .B1(new_n947_), .B2(new_n676_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n953_), .A2(new_n677_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n962_), .B2(new_n331_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1350gat));
  NAND4_X1  g764(.A1(new_n953_), .A2(new_n330_), .A3(new_n332_), .A4(new_n674_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n953_), .A2(new_n715_), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n967_), .A2(KEYINPUT127), .A3(G190gat), .ZN(new_n968_));
  AOI21_X1  g767(.A(KEYINPUT127), .B1(new_n967_), .B2(G190gat), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n966_), .B1(new_n968_), .B2(new_n969_), .ZN(G1351gat));
  AND4_X1   g769(.A1(new_n716_), .A2(new_n945_), .A3(new_n691_), .A4(new_n514_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n971_), .A2(new_n670_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n595_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g774(.A1(new_n971_), .A2(new_n677_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  AND2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  NOR3_X1   g777(.A1(new_n976_), .A2(new_n977_), .A3(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n979_), .B1(new_n976_), .B2(new_n977_), .ZN(G1354gat));
  INV_X1    g779(.A(G218gat), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n971_), .A2(new_n981_), .A3(new_n674_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n971_), .A2(new_n715_), .ZN(new_n983_));
  INV_X1    g782(.A(new_n983_), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n982_), .B1(new_n984_), .B2(new_n981_), .ZN(G1355gat));
endmodule


