//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_;
  AOI21_X1  g000(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT88), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT87), .ZN(new_n204_));
  INV_X1    g003(.A(G141gat), .ZN(new_n205_));
  INV_X1    g004(.A(G148gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  AOI22_X1  g007(.A1(KEYINPUT3), .A2(new_n207_), .B1(new_n208_), .B2(KEYINPUT2), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n203_), .B(new_n209_), .C1(KEYINPUT3), .C2(new_n207_), .ZN(new_n210_));
  INV_X1    g009(.A(G155gat), .ZN(new_n211_));
  INV_X1    g010(.A(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT86), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n210_), .B(new_n214_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n211_), .B2(new_n212_), .ZN(new_n216_));
  OR3_X1    g015(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT1), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n205_), .A2(new_n206_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT28), .ZN(new_n225_));
  INV_X1    g024(.A(G228gat), .ZN(new_n226_));
  INV_X1    g025(.A(G233gat), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n226_), .A2(new_n227_), .A3(KEYINPUT90), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n225_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(G197gat), .B(G204gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT89), .B1(new_n232_), .B2(KEYINPUT21), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n236_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT89), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n235_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n243_));
  INV_X1    g042(.A(G78gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT90), .B1(new_n226_), .B2(new_n227_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n231_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n245_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G78gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G106gat), .A3(new_n246_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G22gat), .B(G50gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n230_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n249_), .A2(new_n252_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n253_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n229_), .A3(new_n255_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT96), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT25), .B(G183gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT77), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT24), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  MUX2_X1   g071(.A(new_n271_), .B(KEYINPUT24), .S(new_n272_), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n268_), .A2(KEYINPUT23), .ZN(new_n275_));
  MUX2_X1   g074(.A(new_n275_), .B(new_n269_), .S(KEYINPUT80), .Z(new_n276_));
  OR2_X1    g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n270_), .ZN(new_n279_));
  AND2_X1   g078(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n280_));
  NOR2_X1   g079(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n281_));
  OAI21_X1  g080(.A(G169gat), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT79), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT22), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(new_n285_), .B2(G169gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n274_), .B1(new_n279_), .B2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(new_n242_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT19), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G169gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n284_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n269_), .A2(new_n277_), .B1(G169gat), .B2(G176gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n273_), .A2(new_n266_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n295_), .A2(new_n296_), .B1(new_n297_), .B2(new_n276_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT20), .B1(new_n298_), .B2(new_n241_), .ZN(new_n299_));
  OR3_X1    g098(.A1(new_n289_), .A2(new_n291_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n288_), .A2(new_n242_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT20), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n298_), .B2(new_n241_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n291_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G8gat), .B(G36gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G64gat), .B(G92gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT27), .ZN(new_n314_));
  INV_X1    g113(.A(new_n291_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n301_), .A2(new_n303_), .A3(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT92), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n291_), .B1(new_n289_), .B2(new_n299_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(KEYINPUT92), .A3(new_n316_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n312_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n263_), .B1(new_n314_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT27), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n319_), .A3(new_n312_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n324_), .B2(new_n320_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n319_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n311_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n327_), .A2(KEYINPUT96), .A3(KEYINPUT27), .A4(new_n313_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n321_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n262_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G15gat), .B(G43gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT82), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G71gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G99gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT83), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n288_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n337_), .A2(new_n340_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n331_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT85), .A3(new_n341_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT84), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT31), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n344_), .A2(new_n346_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n331_), .B(new_n356_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT94), .ZN(new_n360_));
  INV_X1    g159(.A(new_n353_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n222_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n215_), .A2(new_n221_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n353_), .B1(new_n363_), .B2(KEYINPUT94), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n359_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n222_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n364_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n366_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G1gat), .B(G29gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G57gat), .B(G85gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n369_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n371_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n368_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n358_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n330_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n381_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n258_), .A2(new_n261_), .A3(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n321_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n369_), .A2(KEYINPUT33), .A3(new_n371_), .A4(new_n377_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n366_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n365_), .A2(new_n391_), .A3(new_n367_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n370_), .A2(new_n391_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n376_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n327_), .B(new_n323_), .C1(new_n392_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n311_), .A2(KEYINPUT32), .ZN(new_n396_));
  MUX2_X1   g195(.A(new_n306_), .B(new_n326_), .S(new_n396_), .Z(new_n397_));
  OAI22_X1  g196(.A1(new_n390_), .A2(new_n395_), .B1(new_n384_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n258_), .A2(new_n261_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n385_), .A2(new_n386_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n358_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n383_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G29gat), .B(G36gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G43gat), .B(G50gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT73), .B(G15gat), .ZN(new_n411_));
  INV_X1    g210(.A(G22gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT74), .B(G8gat), .Z(new_n414_));
  INV_X1    g213(.A(G1gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT14), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G1gat), .B(G8gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n413_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n410_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT15), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n409_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n407_), .A2(KEYINPUT15), .A3(new_n408_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n421_), .A3(new_n420_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G229gat), .A2(G233gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n423_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n420_), .A2(new_n410_), .A3(new_n421_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n433_), .B2(new_n422_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G113gat), .B(G141gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT76), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G169gat), .B(G197gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n430_), .A2(new_n434_), .A3(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G230gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT64), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G99gat), .A2(G106gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI22_X1  g247(.A1(KEYINPUT70), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(KEYINPUT6), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(KEYINPUT69), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n451_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(KEYINPUT69), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(KEYINPUT6), .ZN(new_n458_));
  AND2_X1   g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n450_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G85gat), .B(G92gat), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT8), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n459_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n449_), .B(new_n448_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n462_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT10), .B(G99gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT65), .B(G106gat), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n456_), .A2(new_n460_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT68), .ZN(new_n474_));
  OR2_X1    g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(KEYINPUT67), .A2(G85gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(KEYINPUT67), .A2(G85gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(G92gat), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT66), .B(KEYINPUT9), .ZN(new_n481_));
  AOI211_X1 g280(.A(new_n474_), .B(new_n477_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n477_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT68), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n473_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G57gat), .B(G64gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G71gat), .B(G78gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT11), .ZN(new_n489_));
  INV_X1    g288(.A(new_n488_), .ZN(new_n490_));
  INV_X1    g289(.A(G64gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G57gat), .ZN(new_n492_));
  INV_X1    g291(.A(G57gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G64gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n494_), .A3(KEYINPUT11), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n487_), .A2(KEYINPUT11), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n489_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n470_), .A2(new_n486_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n470_), .B2(new_n486_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n445_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT68), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n504_), .A2(new_n473_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n487_), .A2(KEYINPUT11), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n495_), .A3(new_n490_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n508_), .B2(new_n489_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n506_), .B(new_n489_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT12), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  OAI22_X1  g311(.A1(new_n501_), .A2(KEYINPUT12), .B1(new_n505_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n445_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n502_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT5), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G176gat), .B(G204gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n502_), .B(new_n522_), .C1(new_n513_), .C2(new_n515_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT13), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n521_), .A2(KEYINPUT13), .A3(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n420_), .A2(new_n421_), .ZN(new_n530_));
  AND2_X1   g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n498_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT16), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT17), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n534_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n509_), .A2(new_n511_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n532_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n532_), .A2(new_n542_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT75), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT75), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n556_), .A2(KEYINPUT36), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n470_), .A2(new_n409_), .A3(new_n486_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n425_), .A2(new_n426_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n470_), .B2(new_n486_), .ZN(new_n563_));
  OAI211_X1 g362(.A(KEYINPUT35), .B(new_n560_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n468_), .B1(new_n467_), .B2(new_n462_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n461_), .A2(KEYINPUT8), .A3(new_n463_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n486_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n427_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n470_), .A2(new_n409_), .A3(new_n486_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n556_), .A2(KEYINPUT36), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n564_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n564_), .B2(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n558_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT37), .B1(new_n574_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n564_), .A2(new_n572_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n564_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n583_), .B2(KEYINPUT72), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n558_), .A3(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n579_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n553_), .A2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n402_), .A2(new_n443_), .A3(new_n529_), .A4(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT97), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT97), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n415_), .A3(new_n381_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n402_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n576_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n443_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n528_), .A2(new_n599_), .A3(new_n548_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n384_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n594_), .A2(new_n595_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n596_), .A2(new_n603_), .A3(new_n604_), .ZN(G1324gat));
  XNOR2_X1  g404(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n606_));
  INV_X1    g405(.A(new_n576_), .ZN(new_n607_));
  AND4_X1   g406(.A1(new_n329_), .A2(new_n402_), .A3(new_n607_), .A4(new_n600_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(G8gat), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n608_), .A2(new_n609_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT39), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AND4_X1   g412(.A1(KEYINPUT39), .A2(new_n612_), .A3(G8gat), .A4(new_n610_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n329_), .A2(new_n414_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n591_), .A2(new_n592_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT98), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n591_), .A2(new_n619_), .A3(new_n592_), .A4(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n606_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(KEYINPUT39), .A3(new_n612_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n612_), .A2(G8gat), .A3(new_n610_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AND4_X1   g425(.A1(new_n621_), .A2(new_n623_), .A3(new_n626_), .A4(new_n606_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n622_), .A2(new_n627_), .ZN(G1325gat));
  OAI21_X1  g427(.A(G15gat), .B1(new_n602_), .B2(new_n358_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n630_), .ZN(new_n632_));
  INV_X1    g431(.A(G15gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n593_), .A2(new_n633_), .A3(new_n401_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n632_), .A3(new_n634_), .ZN(G1326gat));
  AOI21_X1  g434(.A(new_n412_), .B1(new_n601_), .B2(new_n262_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT42), .Z(new_n637_));
  NOR2_X1   g436(.A1(new_n399_), .A2(G22gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT102), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n593_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(G1327gat));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n579_), .A2(new_n587_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT103), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n385_), .A2(new_n386_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n398_), .A2(new_n399_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n401_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NOR4_X1   g446(.A1(new_n262_), .A2(new_n358_), .A3(new_n329_), .A4(new_n381_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n643_), .A2(KEYINPUT43), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n649_), .A2(KEYINPUT43), .B1(new_n402_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n528_), .A2(new_n599_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n553_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n642_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n402_), .A2(new_n650_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n402_), .B2(new_n644_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n655_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n384_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n553_), .A2(new_n576_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n528_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n402_), .A2(new_n443_), .A3(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n384_), .A2(G29gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT104), .ZN(G1328gat));
  NOR2_X1   g466(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n386_), .A2(G36gat), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n664_), .A2(KEYINPUT45), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT45), .B1(new_n664_), .B2(new_n669_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n654_), .A2(new_n329_), .A3(new_n659_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT105), .B1(new_n673_), .B2(G36gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT107), .Z(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n672_), .B(new_n678_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1329gat));
  NAND2_X1  g481(.A1(new_n401_), .A2(G43gat), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n664_), .A2(new_n358_), .ZN(new_n684_));
  OAI22_X1  g483(.A1(new_n660_), .A2(new_n683_), .B1(G43gat), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g485(.A(G50gat), .B1(new_n660_), .B2(new_n399_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n399_), .A2(G50gat), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT108), .Z(new_n689_));
  OAI21_X1  g488(.A(new_n687_), .B1(new_n664_), .B2(new_n689_), .ZN(G1331gat));
  NAND2_X1  g489(.A1(new_n589_), .A2(new_n528_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT109), .Z(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n597_), .A3(new_n443_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n493_), .A3(new_n381_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n549_), .A2(new_n599_), .A3(new_n551_), .ZN(new_n695_));
  NOR4_X1   g494(.A1(new_n597_), .A2(new_n529_), .A3(new_n576_), .A4(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(new_n381_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n697_), .B2(new_n493_), .ZN(G1332gat));
  AOI21_X1  g497(.A(new_n491_), .B1(new_n696_), .B2(new_n329_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n329_), .A2(new_n491_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT111), .Z(new_n703_));
  NAND2_X1  g502(.A1(new_n693_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1333gat));
  INV_X1    g504(.A(G71gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n696_), .B2(new_n401_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT49), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n693_), .A2(new_n706_), .A3(new_n401_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1334gat));
  AOI21_X1  g509(.A(new_n244_), .B1(new_n696_), .B2(new_n262_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT50), .Z(new_n712_));
  NOR2_X1   g511(.A1(new_n399_), .A2(G78gat), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT112), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n693_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1335gat));
  INV_X1    g515(.A(new_n651_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n552_), .A2(new_n529_), .A3(new_n443_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n478_), .A2(new_n479_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n719_), .A2(new_n384_), .A3(new_n720_), .ZN(new_n721_));
  NOR4_X1   g520(.A1(new_n597_), .A2(new_n443_), .A3(new_n529_), .A4(new_n662_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n381_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1336gat));
  OAI21_X1  g523(.A(G92gat), .B1(new_n719_), .B2(new_n386_), .ZN(new_n725_));
  INV_X1    g524(.A(G92gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n726_), .A3(new_n329_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1337gat));
  NOR2_X1   g527(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n729_));
  OAI21_X1  g528(.A(G99gat), .B1(new_n719_), .B2(new_n358_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n722_), .A2(new_n401_), .A3(new_n471_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n732_), .B(new_n733_), .Z(G1338gat));
  NAND3_X1  g533(.A1(new_n722_), .A2(new_n262_), .A3(new_n472_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n717_), .A2(new_n262_), .A3(new_n718_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G106gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g540(.A(KEYINPUT122), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n695_), .A2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n695_), .A2(new_n743_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n528_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n643_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n643_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT54), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n746_), .A2(KEYINPUT115), .A3(new_n747_), .A4(new_n643_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n750_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n548_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n443_), .A2(new_n523_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT12), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n498_), .A2(KEYINPUT71), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n510_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n567_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n499_), .C1(KEYINPUT12), .C2(new_n501_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n445_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n505_), .B2(new_n498_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n445_), .B1(new_n505_), .B2(new_n498_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(KEYINPUT55), .A4(new_n766_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n520_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n520_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n423_), .A2(new_n428_), .A3(new_n431_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n429_), .B1(new_n433_), .B2(new_n422_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n440_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n442_), .A2(new_n780_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n760_), .A2(new_n777_), .B1(new_n524_), .B2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n756_), .B(new_n757_), .C1(new_n782_), .C2(new_n576_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n756_), .A2(new_n757_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n760_), .A2(new_n777_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n524_), .A2(new_n781_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n607_), .B(new_n784_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n781_), .A2(new_n523_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n520_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n520_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT119), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n790_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n801_), .B(new_n643_), .C1(new_n795_), .C2(new_n794_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n794_), .A2(new_n795_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT118), .B1(new_n803_), .B2(new_n588_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n588_), .B1(new_n797_), .B2(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n801_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(KEYINPUT118), .A3(new_n588_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT120), .B1(new_n811_), .B2(new_n800_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n789_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n755_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n805_), .A2(new_n806_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(KEYINPUT120), .A3(new_n800_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n788_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT121), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n754_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n330_), .A2(new_n381_), .A3(new_n401_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n742_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n750_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n548_), .B1(new_n818_), .B2(KEYINPUT121), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n814_), .B(new_n788_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n821_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT122), .A3(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n822_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(G113gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n443_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n789_), .A2(new_n805_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n553_), .ZN(new_n833_));
  AOI211_X1 g632(.A(KEYINPUT59), .B(new_n821_), .C1(new_n833_), .C2(new_n823_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n826_), .A2(new_n827_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(KEYINPUT59), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(new_n443_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n831_), .B1(new_n830_), .B2(new_n837_), .ZN(G1340gat));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n529_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n829_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n839_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n836_), .A2(new_n528_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n839_), .B2(new_n842_), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n829_), .A2(new_n844_), .A3(new_n552_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n836_), .A2(new_n755_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n844_), .B2(new_n846_), .ZN(G1342gat));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n836_), .B2(new_n588_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n607_), .A2(G134gat), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n822_), .A2(new_n828_), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n848_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n822_), .A2(new_n828_), .A3(new_n851_), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n643_), .B(new_n834_), .C1(new_n835_), .C2(KEYINPUT59), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT123), .B(new_n854_), .C1(new_n855_), .C2(new_n849_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1343gat));
  NOR4_X1   g656(.A1(new_n401_), .A2(new_n399_), .A3(new_n329_), .A4(new_n384_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n826_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n599_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n205_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n529_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n206_), .ZN(G1345gat));
  AND2_X1   g662(.A1(new_n826_), .A2(new_n858_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(KEYINPUT124), .A3(new_n552_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n859_), .B2(new_n553_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT125), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n868_), .B(new_n871_), .ZN(G1346gat));
  AOI21_X1  g671(.A(G162gat), .B1(new_n864_), .B2(new_n576_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n644_), .A2(G162gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n864_), .B2(new_n874_), .ZN(G1347gat));
  NAND2_X1  g674(.A1(new_n382_), .A2(new_n329_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n552_), .B1(new_n789_), .B2(new_n805_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n399_), .B(new_n877_), .C1(new_n754_), .C2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879_), .B2(new_n599_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT62), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n879_), .B(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n443_), .A3(new_n294_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n884_), .ZN(G1348gat));
  XNOR2_X1  g684(.A(new_n879_), .B(KEYINPUT126), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n284_), .B1(new_n886_), .B2(new_n529_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n826_), .A2(new_n399_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n877_), .A2(G176gat), .A3(new_n528_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n887_), .B(new_n888_), .C1(new_n889_), .C2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G176gat), .B1(new_n883_), .B2(new_n528_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n890_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT127), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(G1349gat));
  NOR3_X1   g694(.A1(new_n886_), .A2(new_n264_), .A3(new_n548_), .ZN(new_n896_));
  INV_X1    g695(.A(G183gat), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n826_), .A2(new_n399_), .A3(new_n552_), .A4(new_n877_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n886_), .B2(new_n643_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n883_), .A2(new_n265_), .A3(new_n576_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1351gat));
  AND4_X1   g701(.A1(new_n385_), .A2(new_n826_), .A3(new_n329_), .A4(new_n358_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n443_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n528_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n755_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT63), .B(G211gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n908_), .B2(new_n911_), .ZN(G1354gat));
  INV_X1    g711(.A(G218gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n903_), .A2(new_n913_), .A3(new_n576_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n903_), .A2(new_n588_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n913_), .ZN(G1355gat));
endmodule


