//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT21), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT21), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT88), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n214_), .A2(KEYINPUT3), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n216_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT2), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n217_), .B(new_n219_), .C1(new_n223_), .C2(KEYINPUT90), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(KEYINPUT90), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n213_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT91), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(KEYINPUT91), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n212_), .B(KEYINPUT1), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n211_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n218_), .A2(new_n220_), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n227_), .A2(new_n228_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n209_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G228gat), .ZN(new_n235_));
  INV_X1    g034(.A(G233gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  OAI221_X1 g037(.A(new_n209_), .B1(new_n235_), .B2(new_n236_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G78gat), .B(G106gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT92), .Z(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(KEYINPUT93), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G22gat), .B(G50gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT28), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n230_), .A2(new_n231_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n226_), .A2(KEYINPUT91), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n226_), .A2(KEYINPUT91), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n252_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n246_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n232_), .A2(new_n247_), .A3(new_n233_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT28), .B1(new_n252_), .B2(KEYINPUT29), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n245_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n244_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT93), .B1(new_n240_), .B2(new_n243_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT94), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n259_), .A2(new_n257_), .A3(new_n254_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT94), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .A4(new_n244_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n240_), .A2(new_n243_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n268_), .A2(new_n259_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(new_n258_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT23), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT84), .B(KEYINPUT23), .Z(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(new_n273_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(G183gat), .B2(G190gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT22), .B(G169gat), .ZN(new_n278_));
  INV_X1    g077(.A(G176gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT83), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n282_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT25), .B(G183gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G190gat), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n288_), .B2(new_n287_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT85), .B1(new_n273_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n275_), .A2(new_n272_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n273_), .A2(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n297_), .B1(new_n300_), .B2(KEYINPUT85), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n284_), .B1(new_n295_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT86), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT86), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n284_), .B(new_n304_), .C1(new_n295_), .C2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G71gat), .B(G99gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G43gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G127gat), .B(G134gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT87), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G113gat), .B(G120gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n309_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G227gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(G15gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT30), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT31), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n315_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n252_), .A2(new_n314_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n313_), .B(new_n249_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(KEYINPUT4), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n252_), .A2(new_n327_), .A3(new_n314_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G1gat), .B(G29gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT97), .B(G85gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n329_), .A2(new_n330_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n209_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n289_), .A2(new_n281_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n293_), .B1(new_n288_), .B2(new_n285_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n276_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n301_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n283_), .B(KEYINPUT96), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n346_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n350_), .B2(new_n209_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n343_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n350_), .B2(new_n209_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n303_), .A2(new_n342_), .A3(new_n305_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n356_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT18), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n343_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n361_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n359_), .A2(new_n360_), .ZN(new_n374_));
  MUX2_X1   g173(.A(new_n374_), .B(new_n352_), .S(new_n355_), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n366_), .B(KEYINPUT100), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT27), .B(new_n367_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n377_), .ZN(new_n378_));
  NOR4_X1   g177(.A1(new_n271_), .A2(new_n321_), .A3(new_n341_), .A4(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n271_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n337_), .A2(KEYINPUT98), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT33), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n324_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n322_), .A2(new_n323_), .A3(new_n326_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n335_), .A3(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n367_), .A2(new_n385_), .A3(new_n370_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n337_), .A2(KEYINPUT98), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT99), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT99), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n386_), .A3(new_n391_), .A4(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n357_), .A2(new_n362_), .A3(new_n393_), .ZN(new_n394_));
  OAI221_X1 g193(.A(new_n394_), .B1(new_n375_), .B2(new_n393_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n380_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n378_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n340_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n379_), .B1(new_n400_), .B2(new_n321_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G29gat), .B(G36gat), .Z(new_n402_));
  XOR2_X1   g201(.A(G43gat), .B(G50gat), .Z(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT15), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT75), .B(G8gat), .ZN(new_n406_));
  INV_X1    g205(.A(G1gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT14), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G15gat), .B(G22gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G8gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n405_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n404_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n415_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G229gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n415_), .B(new_n404_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT79), .Z(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n425_), .B2(new_n420_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G113gat), .B(G141gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT80), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G169gat), .B(G197gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n428_), .B(new_n429_), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n423_), .B(new_n430_), .C1(new_n425_), .C2(new_n420_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n426_), .A2(KEYINPUT81), .A3(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT68), .B(G71gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G78gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G57gat), .B(G64gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT11), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n440_), .A2(KEYINPUT11), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G78gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n438_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n441_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n449_));
  AND2_X1   g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G85gat), .A2(G92gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G99gat), .A3(G106gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n452_), .B1(new_n457_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n452_), .A2(KEYINPUT67), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n454_), .A2(new_n456_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n462_), .A3(new_n461_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(new_n466_), .A3(new_n452_), .A4(new_n465_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT10), .B(G99gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n469_), .B1(new_n473_), .B2(G106gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n451_), .B1(new_n450_), .B2(KEYINPUT9), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n476_), .A2(KEYINPUT64), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT64), .B1(new_n476_), .B2(new_n477_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n475_), .B(KEYINPUT65), .C1(new_n478_), .C2(new_n479_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n474_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n472_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AOI211_X1 g285(.A(KEYINPUT66), .B(new_n474_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n448_), .B(new_n449_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n448_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n474_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n479_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n476_), .A2(KEYINPUT64), .A3(new_n477_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT65), .B1(new_n493_), .B2(new_n475_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n483_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n490_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n496_), .A2(KEYINPUT66), .B1(new_n468_), .B2(new_n471_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n484_), .A2(new_n485_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n489_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT69), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT12), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n488_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n486_), .A2(new_n448_), .A3(new_n487_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT70), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G230gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n496_), .A2(KEYINPUT66), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n489_), .A2(new_n508_), .A3(new_n498_), .A4(new_n472_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT70), .B1(new_n509_), .B2(new_n505_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n502_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n499_), .A2(new_n503_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G120gat), .B(G148gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G176gat), .B(G204gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n511_), .B(new_n518_), .C1(new_n505_), .C2(new_n512_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT13), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT13), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT72), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n486_), .A2(new_n487_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(new_n405_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT34), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n417_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n531_), .A2(new_n532_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT73), .ZN(new_n541_));
  XOR2_X1   g340(.A(G134gat), .B(G162gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT36), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n537_), .A2(new_n546_), .A3(new_n543_), .A4(new_n538_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n544_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT37), .B1(new_n550_), .B2(KEYINPUT74), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n548_), .B(new_n551_), .Z(new_n552_));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n415_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n489_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G183gat), .B(G211gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n555_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT77), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n560_), .A2(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT78), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n562_), .B(new_n565_), .C1(new_n555_), .C2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n555_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n552_), .A2(new_n570_), .ZN(new_n571_));
  NOR4_X1   g370(.A1(new_n401_), .A2(new_n437_), .A3(new_n526_), .A4(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(KEYINPUT101), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT101), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n407_), .A3(new_n341_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n548_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n401_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n525_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n570_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n582_), .A2(new_n437_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n340_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n575_), .A2(new_n407_), .A3(new_n341_), .A4(new_n577_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n579_), .A2(new_n586_), .A3(new_n587_), .ZN(G1324gat));
  NAND4_X1  g387(.A1(new_n573_), .A2(new_n378_), .A3(new_n406_), .A4(new_n574_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n378_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT39), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n591_), .A2(new_n592_), .A3(G8gat), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n591_), .B2(G8gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n589_), .B(KEYINPUT40), .C1(new_n593_), .C2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(G1325gat));
  INV_X1    g398(.A(new_n321_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n590_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G15gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT103), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n604_), .A3(G15gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT41), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(KEYINPUT41), .A3(new_n605_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n575_), .A2(new_n317_), .A3(new_n600_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(G1326gat));
  INV_X1    g410(.A(G22gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n575_), .A2(new_n612_), .A3(new_n271_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G22gat), .B1(new_n585_), .B2(new_n380_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(G1327gat));
  INV_X1    g415(.A(KEYINPUT43), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT104), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n548_), .B(new_n551_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n600_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n620_), .B2(new_n379_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(KEYINPUT104), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n618_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n271_), .A2(new_n378_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n340_), .A3(new_n600_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n380_), .A2(new_n396_), .B1(new_n398_), .B2(new_n340_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n625_), .B(new_n627_), .C1(new_n628_), .C2(new_n600_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n617_), .A2(KEYINPUT105), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n629_), .B(new_n619_), .C1(new_n401_), .C2(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n582_), .A2(new_n437_), .A3(new_n570_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n624_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n624_), .A2(new_n631_), .A3(KEYINPUT44), .A4(new_n632_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n341_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(G29gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n627_), .B1(new_n628_), .B2(new_n600_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n437_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n583_), .A2(new_n580_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n582_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n340_), .A2(G29gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT107), .Z(new_n645_));
  OAI21_X1  g444(.A(new_n638_), .B1(new_n643_), .B2(new_n645_), .ZN(G1328gat));
  NAND3_X1  g445(.A1(new_n635_), .A2(new_n378_), .A3(new_n636_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G36gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n378_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n643_), .A2(G36gat), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(new_n652_), .A3(KEYINPUT46), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1329gat));
  NAND4_X1  g456(.A1(new_n635_), .A2(G43gat), .A3(new_n600_), .A4(new_n636_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n643_), .A2(new_n321_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(G43gat), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g460(.A1(new_n635_), .A2(G50gat), .A3(new_n271_), .A4(new_n636_), .ZN(new_n662_));
  INV_X1    g461(.A(G50gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n643_), .B2(new_n380_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1331gat));
  INV_X1    g464(.A(KEYINPUT109), .ZN(new_n666_));
  INV_X1    g465(.A(new_n526_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n437_), .A2(new_n570_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n581_), .A2(new_n666_), .A3(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n639_), .A3(new_n548_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT109), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n670_), .A2(new_n672_), .A3(G57gat), .A4(new_n341_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n673_), .A2(new_n674_), .ZN(new_n676_));
  NOR4_X1   g475(.A1(new_n401_), .A2(new_n640_), .A3(new_n525_), .A4(new_n571_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G57gat), .B1(new_n677_), .B2(new_n341_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n675_), .A2(new_n676_), .A3(new_n678_), .ZN(G1332gat));
  INV_X1    g478(.A(G64gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n680_), .A3(new_n378_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n670_), .A2(new_n672_), .A3(new_n378_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT48), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G64gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G64gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n677_), .A2(new_n687_), .A3(new_n600_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n670_), .A2(new_n672_), .A3(new_n600_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT49), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(G71gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n689_), .B2(G71gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(G1334gat));
  NAND3_X1  g492(.A1(new_n677_), .A2(new_n445_), .A3(new_n271_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n670_), .A2(new_n672_), .A3(new_n271_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT50), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(G78gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G78gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(G1335gat));
  NOR3_X1   g500(.A1(new_n525_), .A2(new_n640_), .A3(new_n570_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n624_), .A2(new_n631_), .A3(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n340_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n401_), .A2(new_n640_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n667_), .A2(new_n641_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(KEYINPUT112), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT112), .B1(new_n705_), .B2(new_n706_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G85gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n341_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n704_), .B1(new_n709_), .B2(new_n711_), .ZN(G1336gat));
  OAI21_X1  g511(.A(G92gat), .B1(new_n703_), .B2(new_n649_), .ZN(new_n713_));
  INV_X1    g512(.A(G92gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n378_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n709_), .B2(new_n715_), .ZN(G1337gat));
  OAI21_X1  g515(.A(G99gat), .B1(new_n703_), .B2(new_n321_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n321_), .A2(new_n473_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT114), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(KEYINPUT114), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n717_), .A2(new_n719_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT51), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n723_), .A3(new_n725_), .ZN(G1338gat));
  NAND4_X1  g525(.A1(new_n624_), .A2(new_n631_), .A3(new_n271_), .A4(new_n702_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G106gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G106gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n271_), .A2(new_n460_), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n729_), .A2(new_n730_), .B1(new_n709_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n732_), .B(new_n734_), .ZN(G1339gat));
  NOR2_X1   g534(.A1(new_n419_), .A2(new_n420_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n430_), .B1(new_n416_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n425_), .B2(new_n421_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n434_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n522_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n522_), .B2(new_n739_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n435_), .A2(new_n436_), .A3(new_n521_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n502_), .A2(new_n509_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n506_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n502_), .B(new_n749_), .C1(new_n507_), .C2(new_n510_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n504_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n509_), .A2(KEYINPUT70), .A3(new_n505_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n749_), .B1(new_n754_), .B2(new_n502_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n746_), .B(new_n748_), .C1(new_n751_), .C2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n519_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n511_), .A2(KEYINPUT55), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n750_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n746_), .B1(new_n759_), .B2(new_n748_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n745_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n748_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT117), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(KEYINPUT56), .A3(new_n519_), .A4(new_n756_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n744_), .B1(new_n761_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n743_), .B1(new_n765_), .B2(KEYINPUT118), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n767_), .B(new_n744_), .C1(new_n761_), .C2(new_n764_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n548_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT57), .B(new_n548_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n739_), .A2(new_n521_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n761_), .B2(new_n764_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(KEYINPUT58), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(KEYINPUT58), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n619_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n771_), .A2(new_n772_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n583_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT122), .ZN(new_n780_));
  INV_X1    g579(.A(new_n668_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n525_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n552_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT116), .B1(new_n781_), .B2(new_n525_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n784_), .A2(KEYINPUT54), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n668_), .B1(new_n524_), .B2(new_n523_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n619_), .B1(new_n788_), .B2(KEYINPUT116), .ZN(new_n789_));
  INV_X1    g588(.A(new_n785_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n786_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n778_), .A2(new_n794_), .A3(new_n583_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n780_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n626_), .A2(new_n341_), .A3(new_n600_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT121), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802_));
  INV_X1    g601(.A(new_n776_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n619_), .B1(new_n774_), .B2(KEYINPUT58), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n775_), .A2(KEYINPUT120), .A3(new_n619_), .A4(new_n776_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n771_), .A2(new_n772_), .A3(new_n805_), .A4(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n583_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n801_), .B1(new_n808_), .B2(new_n793_), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT121), .B(new_n792_), .C1(new_n807_), .C2(new_n583_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n798_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n640_), .B(new_n800_), .C1(new_n811_), .C2(new_n797_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G113gat), .ZN(new_n813_));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n814_), .A3(new_n640_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1340gat));
  OAI211_X1 g615(.A(new_n526_), .B(new_n800_), .C1(new_n811_), .C2(new_n797_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G120gat), .ZN(new_n818_));
  INV_X1    g617(.A(new_n809_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n810_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n525_), .A2(KEYINPUT60), .ZN(new_n821_));
  MUX2_X1   g620(.A(new_n821_), .B(KEYINPUT60), .S(G120gat), .Z(new_n822_));
  NAND4_X1  g621(.A1(new_n819_), .A2(new_n820_), .A3(new_n799_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT123), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n811_), .A2(new_n825_), .A3(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n818_), .A2(new_n827_), .ZN(G1341gat));
  OAI211_X1 g627(.A(new_n570_), .B(new_n800_), .C1(new_n811_), .C2(new_n797_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G127gat), .ZN(new_n830_));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n811_), .A2(new_n831_), .A3(new_n570_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1342gat));
  OAI211_X1 g632(.A(new_n619_), .B(new_n800_), .C1(new_n811_), .C2(new_n797_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G134gat), .ZN(new_n835_));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n811_), .A2(new_n836_), .A3(new_n580_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1343gat));
  NOR2_X1   g637(.A1(new_n809_), .A2(new_n810_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n398_), .A2(new_n341_), .A3(new_n321_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n640_), .A3(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n526_), .A3(new_n840_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT124), .B(G148gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1345gat));
  NAND3_X1  g644(.A1(new_n839_), .A2(new_n570_), .A3(new_n840_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  NAND3_X1  g647(.A1(new_n839_), .A2(new_n619_), .A3(new_n840_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G162gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n548_), .A2(G162gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n839_), .A2(new_n840_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1347gat));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n649_), .A2(new_n341_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n600_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n271_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n796_), .A2(new_n640_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G169gat), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT125), .B(new_n854_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n861_), .B2(KEYINPUT62), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n796_), .A2(new_n857_), .ZN(new_n863_));
  OAI221_X1 g662(.A(new_n862_), .B1(new_n861_), .B2(KEYINPUT62), .C1(new_n863_), .C2(new_n437_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n858_), .A2(new_n278_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n860_), .A2(new_n864_), .A3(new_n865_), .ZN(G1348gat));
  INV_X1    g665(.A(new_n863_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G176gat), .B1(new_n867_), .B2(new_n582_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n809_), .A2(new_n810_), .A3(new_n271_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n667_), .A2(new_n279_), .A3(new_n856_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  NOR3_X1   g670(.A1(new_n863_), .A2(new_n291_), .A3(new_n583_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n869_), .A2(new_n600_), .A3(new_n570_), .A4(new_n855_), .ZN(new_n873_));
  INV_X1    g672(.A(G183gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1350gat));
  OAI21_X1  g674(.A(G190gat), .B1(new_n863_), .B2(new_n552_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n580_), .A2(new_n292_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n863_), .B2(new_n877_), .ZN(G1351gat));
  NAND3_X1  g677(.A1(new_n271_), .A2(new_n855_), .A3(new_n321_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n839_), .A2(new_n640_), .A3(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g681(.A1(new_n839_), .A2(new_n526_), .A3(new_n880_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g683(.A(KEYINPUT63), .B(G211gat), .Z(new_n885_));
  AND4_X1   g684(.A1(new_n570_), .A2(new_n839_), .A3(new_n880_), .A4(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n839_), .A2(new_n570_), .A3(new_n880_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1354gat));
  NAND2_X1  g688(.A1(new_n619_), .A2(G218gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT127), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n809_), .A2(new_n810_), .A3(new_n879_), .A4(new_n891_), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n809_), .A2(new_n810_), .A3(new_n548_), .A4(new_n879_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  AOI21_X1  g693(.A(G218gat), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n839_), .A2(new_n580_), .A3(new_n880_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n892_), .B1(new_n895_), .B2(new_n897_), .ZN(G1355gat));
endmodule


