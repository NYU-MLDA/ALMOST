//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n584_, new_n585_, new_n586_, new_n587_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G155gat), .B(G162gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT85), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n212_), .A2(new_n215_), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n217_), .C1(G141gat), .C2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G134gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT82), .B(G127gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT91), .B1(new_n219_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(new_n223_), .B2(new_n219_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT91), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n219_), .A2(new_n226_), .A3(new_n223_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n202_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G225gat), .A2(G233gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT92), .Z(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n219_), .A2(new_n202_), .A3(new_n223_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n230_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G1gat), .B(G29gat), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G57gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n235_), .A2(KEYINPUT33), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT33), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT90), .ZN(new_n245_));
  OR3_X1    g044(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT24), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n246_), .A2(KEYINPUT24), .A3(new_n253_), .A4(new_n247_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT88), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT25), .B(G183gat), .Z(new_n257_));
  OAI211_X1 g056(.A(new_n252_), .B(new_n254_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n251_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(G183gat), .B2(G190gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT22), .B(G169gat), .ZN(new_n261_));
  INV_X1    g060(.A(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n253_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(G197gat), .B(G204gat), .Z(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(KEYINPUT21), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(KEYINPUT21), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  OR2_X1    g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT20), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  INV_X1    g072(.A(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT22), .ZN(new_n275_));
  AOI21_X1  g074(.A(G176gat), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  OAI221_X1 g075(.A(new_n260_), .B1(new_n273_), .B2(new_n263_), .C1(new_n274_), .C2(new_n276_), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n248_), .A2(new_n251_), .A3(KEYINPUT79), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT79), .B1(new_n248_), .B2(new_n251_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n257_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n255_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n254_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n283_), .A2(new_n270_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT19), .ZN(new_n286_));
  OR3_X1    g085(.A1(new_n272_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G8gat), .B(G36gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  NAND2_X1  g091(.A1(new_n265_), .A2(new_n270_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n293_), .B(KEYINPUT20), .C1(new_n283_), .C2(new_n270_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n286_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n287_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n287_), .B2(new_n295_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n245_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n242_), .A2(new_n244_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT93), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n228_), .A2(new_n232_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(new_n231_), .ZN(new_n303_));
  NOR4_X1   g102(.A1(new_n228_), .A2(KEYINPUT93), .A3(new_n230_), .A4(new_n232_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n231_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n240_), .B1(new_n306_), .B2(new_n243_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n298_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(KEYINPUT90), .A3(new_n296_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n287_), .A2(new_n295_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(KEYINPUT32), .B2(new_n292_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n235_), .A2(new_n241_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n240_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n294_), .A2(new_n286_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n272_), .A2(KEYINPUT94), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT94), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n271_), .B2(KEYINPUT20), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n317_), .A2(new_n284_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n286_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n316_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(KEYINPUT32), .A3(new_n292_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n270_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G106gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(G78gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n330_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT87), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G22gat), .B(G50gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n336_), .A3(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n336_), .A2(new_n341_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n315_), .A2(new_n323_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n310_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT27), .B1(new_n308_), .B2(new_n296_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n292_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n297_), .B1(new_n322_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n348_), .B2(KEYINPUT27), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n313_), .A2(KEYINPUT95), .A3(new_n314_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT95), .B1(new_n313_), .B2(new_n314_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n342_), .A2(new_n343_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n283_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  INV_X1    g157(.A(G15gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n357_), .A2(new_n361_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n362_), .B2(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n355_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n366_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n365_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT83), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n223_), .B(KEYINPUT31), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n369_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n372_), .A2(KEYINPUT83), .A3(new_n373_), .A4(new_n375_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT84), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT84), .B1(new_n377_), .B2(new_n378_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n345_), .A2(new_n354_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT96), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT96), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n345_), .A2(new_n354_), .A3(new_n381_), .A4(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n353_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n349_), .A2(new_n386_), .A3(KEYINPUT97), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT97), .ZN(new_n388_));
  INV_X1    g187(.A(new_n349_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n388_), .B1(new_n353_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n350_), .A2(new_n351_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n377_), .A2(new_n378_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n383_), .A2(new_n385_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G229gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G15gat), .B(G22gat), .Z(new_n399_));
  NAND2_X1  g198(.A1(G1gat), .A2(G8gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(KEYINPUT14), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT71), .ZN(new_n402_));
  XOR2_X1   g201(.A(G1gat), .B(G8gat), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT71), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n401_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G43gat), .B(G50gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(G29gat), .B(G36gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n404_), .A2(new_n408_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n396_), .B(new_n398_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n404_), .A2(new_n408_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n411_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n411_), .B(KEYINPUT15), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n418_), .B(new_n397_), .C1(new_n416_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n412_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n396_), .B1(new_n422_), .B2(new_n398_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G169gat), .B(G197gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G141gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT77), .B(G113gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n421_), .A2(new_n423_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n398_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT75), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n428_), .A2(new_n424_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n420_), .A4(new_n415_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G57gat), .ZN(new_n435_));
  INV_X1    g234(.A(G64gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G57gat), .A2(G64gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT11), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G71gat), .B(G78gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT11), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n437_), .A2(new_n443_), .A3(new_n438_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n441_), .A3(KEYINPUT11), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  INV_X1    g248(.A(G99gat), .ZN(new_n450_));
  INV_X1    g249(.A(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n452_), .A2(new_n455_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G85gat), .B(G92gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n458_), .A2(new_n460_), .A3(new_n461_), .A4(new_n463_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT10), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(G99gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n450_), .A2(KEYINPUT10), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT64), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n450_), .A2(KEYINPUT10), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(G99gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT64), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(G106gat), .B1(new_n471_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G85gat), .A3(G92gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n455_), .B(new_n456_), .C1(new_n459_), .C2(new_n477_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n476_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n448_), .B1(new_n467_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483_));
  INV_X1    g282(.A(new_n475_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n474_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n451_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n480_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n478_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n465_), .A3(new_n466_), .A4(new_n447_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n483_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G230gat), .A2(G233gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n490_), .B(new_n492_), .C1(new_n483_), .C2(new_n489_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n482_), .A2(KEYINPUT12), .A3(new_n489_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n448_), .C1(new_n467_), .C2(new_n481_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n492_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT67), .B(G204gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT5), .B(G176gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G120gat), .B(G148gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n505_), .A2(KEYINPUT68), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT68), .B1(new_n505_), .B2(new_n507_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT13), .ZN(new_n510_));
  OR3_X1    g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n510_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n395_), .A2(new_n434_), .A3(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n467_), .A2(new_n481_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n417_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT34), .ZN(new_n518_));
  OAI221_X1 g317(.A(new_n516_), .B1(KEYINPUT35), .B2(new_n518_), .C1(new_n419_), .C2(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT35), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT69), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(new_n522_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n523_), .A2(KEYINPUT70), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT70), .B1(new_n523_), .B2(new_n524_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G190gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT36), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n525_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n524_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT37), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n530_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(KEYINPUT37), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n447_), .B(new_n544_), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n416_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G183gat), .B(G211gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G127gat), .B(G155gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT73), .Z(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n552_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n546_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT74), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n543_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n514_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(G1gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n392_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT38), .ZN(new_n565_));
  INV_X1    g364(.A(new_n538_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(new_n560_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n514_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n568_), .A2(new_n392_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n563_), .B2(new_n569_), .ZN(G1324gat));
  INV_X1    g369(.A(G8gat), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n562_), .A2(new_n571_), .A3(new_n389_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT98), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n568_), .B2(new_n389_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT39), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(G1325gat));
  INV_X1    g377(.A(new_n381_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n359_), .B1(new_n568_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT41), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n562_), .A2(new_n359_), .A3(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(G1326gat));
  INV_X1    g382(.A(G22gat), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n568_), .B2(new_n353_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT42), .Z(new_n586_));
  NAND3_X1  g385(.A1(new_n562_), .A2(new_n584_), .A3(new_n353_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(G1327gat));
  INV_X1    g387(.A(new_n560_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n538_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT101), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n514_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(G29gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n392_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT102), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n392_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n513_), .A2(new_n434_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT43), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n383_), .A2(new_n385_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n391_), .A2(new_n394_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n599_), .B1(new_n602_), .B2(new_n543_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n543_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n395_), .A2(KEYINPUT43), .A3(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n598_), .B(new_n560_), .C1(new_n603_), .C2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n599_), .A3(new_n543_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT43), .B1(new_n395_), .B2(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(new_n598_), .A3(new_n560_), .A4(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n597_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n596_), .B1(new_n614_), .B2(new_n593_), .ZN(G1328gat));
  INV_X1    g414(.A(KEYINPUT46), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n608_), .A2(new_n613_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT103), .B1(new_n617_), .B2(new_n389_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619_));
  AOI211_X1 g418(.A(new_n619_), .B(new_n349_), .C1(new_n608_), .C2(new_n613_), .ZN(new_n620_));
  INV_X1    g419(.A(G36gat), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n618_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n592_), .A2(new_n621_), .A3(new_n389_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT45), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n616_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n618_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n620_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(G36gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(KEYINPUT46), .A3(new_n624_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(G1329gat));
  NAND3_X1  g430(.A1(new_n592_), .A2(new_n364_), .A3(new_n579_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n393_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(new_n364_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g434(.A(G50gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n592_), .A2(new_n636_), .A3(new_n353_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n386_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n636_), .ZN(G1331gat));
  NAND2_X1  g438(.A1(new_n513_), .A2(new_n434_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n395_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(new_n561_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G57gat), .B1(new_n642_), .B2(new_n392_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n641_), .A2(new_n567_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n597_), .A2(new_n435_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(G1332gat));
  AOI21_X1  g445(.A(new_n436_), .B1(new_n644_), .B2(new_n389_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT48), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(new_n436_), .A3(new_n389_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1333gat));
  INV_X1    g449(.A(G71gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n644_), .B2(new_n579_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT49), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n642_), .A2(new_n651_), .A3(new_n579_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1334gat));
  AOI21_X1  g454(.A(new_n328_), .B1(new_n644_), .B2(new_n353_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT50), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n642_), .A2(new_n328_), .A3(new_n353_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1335gat));
  NAND2_X1  g458(.A1(new_n641_), .A2(new_n591_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT104), .ZN(new_n661_));
  AOI21_X1  g460(.A(G85gat), .B1(new_n661_), .B2(new_n392_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n611_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n513_), .A2(new_n434_), .A3(new_n560_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n597_), .A2(new_n237_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n662_), .B1(new_n667_), .B2(new_n668_), .ZN(G1336gat));
  AOI21_X1  g468(.A(G92gat), .B1(new_n661_), .B2(new_n389_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT106), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n389_), .A2(G92gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n667_), .B2(new_n672_), .ZN(G1337gat));
  AOI21_X1  g472(.A(new_n450_), .B1(new_n667_), .B2(new_n579_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT51), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n471_), .A2(new_n475_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n393_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n661_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n675_), .A2(new_n676_), .A3(new_n680_), .A4(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n680_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT51), .B1(new_n683_), .B2(new_n674_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1338gat));
  NAND3_X1  g484(.A1(new_n661_), .A2(new_n451_), .A3(new_n353_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n611_), .A2(new_n353_), .A3(new_n560_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G106gat), .B1(new_n687_), .B2(new_n640_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT52), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT52), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g491(.A1(new_n495_), .A2(new_n497_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n491_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT108), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n495_), .A2(new_n492_), .A3(new_n497_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT55), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n498_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n696_), .A2(KEYINPUT55), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n698_), .B1(new_n693_), .B2(new_n491_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT108), .B(new_n492_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(new_n704_), .A3(new_n506_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT56), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n700_), .A2(new_n704_), .A3(KEYINPUT56), .A4(new_n506_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n434_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n505_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n416_), .A2(new_n419_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n398_), .B1(new_n714_), .B2(new_n414_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n418_), .A2(new_n397_), .A3(new_n412_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n428_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n421_), .A2(new_n423_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n428_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n434_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(KEYINPUT109), .A3(new_n505_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT57), .B1(new_n723_), .B2(new_n538_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT58), .ZN(new_n725_));
  INV_X1    g524(.A(new_n708_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n707_), .A2(KEYINPUT110), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n705_), .A2(new_n728_), .A3(new_n706_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n719_), .A2(new_n505_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n725_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n729_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n728_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n708_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n731_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT58), .A3(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n732_), .A2(new_n543_), .A3(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n724_), .A2(new_n738_), .ZN(new_n739_));
  AND4_X1   g538(.A1(KEYINPUT109), .A2(new_n709_), .A3(new_n710_), .A4(new_n505_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT109), .B1(new_n721_), .B2(new_n505_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n566_), .B1(new_n742_), .B2(new_n720_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT57), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n589_), .B1(new_n739_), .B2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n540_), .A2(new_n434_), .A3(new_n589_), .A4(new_n542_), .ZN(new_n746_));
  OR3_X1    g545(.A1(new_n746_), .A2(new_n513_), .A3(KEYINPUT54), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT54), .B1(new_n746_), .B2(new_n513_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n745_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n391_), .A2(new_n392_), .A3(new_n678_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G113gat), .B1(new_n753_), .B2(new_n710_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT59), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n732_), .A2(new_n543_), .A3(new_n737_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT112), .B(new_n757_), .C1(new_n743_), .C2(KEYINPUT57), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n724_), .B2(new_n738_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n760_), .A3(new_n744_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n750_), .B1(new_n761_), .B2(new_n560_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT111), .B(KEYINPUT59), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n762_), .A2(new_n752_), .A3(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n756_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT113), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n710_), .A2(G113gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n754_), .B1(new_n766_), .B2(new_n767_), .ZN(G1340gat));
  XOR2_X1   g567(.A(KEYINPUT114), .B(G120gat), .Z(new_n769_));
  INV_X1    g568(.A(new_n513_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(KEYINPUT60), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n753_), .B(new_n771_), .C1(KEYINPUT60), .C2(new_n769_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT115), .Z(new_n773_));
  NOR3_X1   g572(.A1(new_n756_), .A2(new_n764_), .A3(new_n770_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n769_), .ZN(G1341gat));
  AOI21_X1  g574(.A(G127gat), .B1(new_n753_), .B2(new_n589_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n589_), .A2(G127gat), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n766_), .B2(new_n778_), .ZN(G1342gat));
  AOI21_X1  g578(.A(G134gat), .B1(new_n753_), .B2(new_n566_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n543_), .A2(G134gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n766_), .B2(new_n781_), .ZN(G1343gat));
  NOR3_X1   g581(.A1(new_n751_), .A2(new_n386_), .A3(new_n579_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n392_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT116), .B1(new_n784_), .B2(new_n389_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n783_), .A2(new_n786_), .A3(new_n392_), .A4(new_n349_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n710_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n513_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT117), .B(G148gat), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(G1345gat));
  INV_X1    g592(.A(G155gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n788_), .A2(new_n794_), .A3(new_n589_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT118), .B(KEYINPUT61), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n794_), .B1(new_n788_), .B2(new_n589_), .ZN(new_n799_));
  OR3_X1    g598(.A1(new_n796_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1346gat));
  INV_X1    g601(.A(G162gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n788_), .A2(new_n803_), .A3(new_n566_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n604_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT119), .ZN(G1347gat));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n392_), .A2(new_n349_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n579_), .A2(new_n810_), .A3(new_n386_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n761_), .A2(new_n560_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n749_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n809_), .B1(new_n813_), .B2(new_n710_), .ZN(new_n814_));
  NOR4_X1   g613(.A1(new_n762_), .A2(KEYINPUT120), .A3(new_n434_), .A4(new_n811_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n274_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n808_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n817_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n812_), .A2(new_n749_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n811_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n710_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n813_), .A2(new_n809_), .A3(new_n710_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(G169gat), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT121), .A3(KEYINPUT62), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n818_), .A2(new_n819_), .A3(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n813_), .B(KEYINPUT122), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n710_), .A3(new_n261_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(KEYINPUT123), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1348gat));
  NAND2_X1  g633(.A1(new_n828_), .A2(new_n513_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n262_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n836_), .A2(KEYINPUT124), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(KEYINPUT124), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n751_), .A2(new_n811_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n770_), .A2(new_n262_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n837_), .A2(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1349gat));
  AOI21_X1  g640(.A(G183gat), .B1(new_n839_), .B2(new_n589_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n589_), .A2(new_n257_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n828_), .B2(new_n844_), .ZN(G1350gat));
  INV_X1    g644(.A(new_n256_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n828_), .A2(new_n846_), .A3(new_n566_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n828_), .A2(new_n543_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G190gat), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n849_), .A2(KEYINPUT125), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(KEYINPUT125), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n847_), .B1(new_n850_), .B2(new_n851_), .ZN(G1351gat));
  NAND2_X1  g651(.A1(new_n783_), .A2(new_n810_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n434_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT126), .B(G197gat), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1352gat));
  NOR2_X1   g655(.A1(new_n853_), .A2(new_n770_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1353gat));
  INV_X1    g658(.A(new_n853_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n589_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  AND2_X1   g661(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n861_), .B2(new_n862_), .ZN(G1354gat));
  INV_X1    g664(.A(G218gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n853_), .A2(new_n866_), .A3(new_n604_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n860_), .A2(new_n566_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n866_), .B2(new_n868_), .ZN(G1355gat));
endmodule


