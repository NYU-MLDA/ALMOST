//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n805_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  MUX2_X1   g005(.A(new_n206_), .B(new_n205_), .S(KEYINPUT82), .Z(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT79), .B(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(G190gat), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT81), .B(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT22), .B1(new_n212_), .B2(KEYINPUT80), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n212_), .A2(KEYINPUT22), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n213_), .C1(new_n214_), .C2(KEYINPUT80), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(KEYINPUT24), .B2(new_n219_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n209_), .B2(KEYINPUT25), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n222_), .B(new_n206_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(G71gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n228_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G15gat), .B(G43gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT83), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT30), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n235_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT85), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G113gat), .B(G120gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT84), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n236_), .A2(KEYINPUT85), .A3(new_n237_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n238_), .A2(new_n243_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G197gat), .B(G204gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n250_), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT89), .Z(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G155gat), .B(G162gat), .Z(new_n260_));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT86), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n269_), .A2(new_n271_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n260_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n267_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT29), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n259_), .A2(KEYINPUT88), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G106gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n278_), .A2(G106gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(G78gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n276_), .A2(KEYINPUT29), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G22gat), .B(G50gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT91), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(KEYINPUT91), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n248_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT20), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT25), .B(G183gat), .Z(new_n302_));
  OAI211_X1 g101(.A(new_n207_), .B(new_n222_), .C1(new_n226_), .C2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n211_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n216_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n301_), .B1(new_n259_), .B2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n259_), .B2(new_n228_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT19), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n259_), .A2(new_n308_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n301_), .B1(new_n259_), .B2(new_n228_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n312_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G8gat), .B(G36gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT93), .ZN(new_n321_));
  XOR2_X1   g120(.A(G64gat), .B(G92gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n327_));
  INV_X1    g126(.A(new_n325_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n318_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n319_), .A2(new_n327_), .A3(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n241_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n276_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n241_), .A2(new_n267_), .A3(new_n275_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n336_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT4), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT95), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n276_), .A3(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n338_), .B1(new_n344_), .B2(new_n337_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT0), .B(G57gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n345_), .A2(KEYINPUT33), .A3(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n337_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n349_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT97), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n336_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(G225gat), .B(G233gat), .C1(new_n339_), .C2(KEYINPUT97), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n354_), .B(new_n355_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n332_), .A2(new_n352_), .A3(new_n353_), .A4(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n345_), .A2(new_n349_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n350_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n325_), .A2(KEYINPUT32), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n318_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n259_), .B1(KEYINPUT98), .B2(new_n308_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(KEYINPUT98), .B2(new_n308_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n316_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n312_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n312_), .B2(new_n310_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n364_), .B1(new_n369_), .B2(new_n363_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n300_), .B1(new_n360_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n330_), .A2(new_n373_), .A3(new_n331_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n328_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(KEYINPUT27), .A3(new_n326_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n246_), .A2(new_n245_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n296_), .B(new_n298_), .C1(new_n379_), .C2(new_n244_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n299_), .A2(new_n247_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n362_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n372_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT75), .B(G1gat), .ZN(new_n384_));
  INV_X1    g183(.A(G8gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT14), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G15gat), .B(G22gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G1gat), .B(G8gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G29gat), .B(G36gat), .Z(new_n393_));
  XOR2_X1   g192(.A(G43gat), .B(G50gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n392_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G229gat), .A2(G233gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT15), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n395_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n392_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n406_), .A3(new_n400_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G113gat), .B(G141gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT78), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G169gat), .B(G197gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n402_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G232gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT35), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G85gat), .B(G92gat), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT65), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT65), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT6), .ZN(new_n428_));
  AND2_X1   g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT7), .ZN(new_n434_));
  AOI211_X1 g233(.A(KEYINPUT8), .B(new_n424_), .C1(new_n432_), .C2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT7), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n433_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439_));
  INV_X1    g238(.A(new_n429_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n427_), .A2(KEYINPUT6), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n425_), .A2(KEYINPUT65), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n438_), .B1(new_n439_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(KEYINPUT67), .A3(new_n444_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n424_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT8), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n436_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT64), .B(G85gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G92gat), .ZN(new_n453_));
  OR3_X1    g252(.A1(new_n452_), .A2(KEYINPUT9), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n423_), .A2(KEYINPUT9), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT10), .B(G99gat), .Z(new_n456_));
  INV_X1    g255(.A(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n454_), .A2(new_n432_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n404_), .B1(new_n450_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n439_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n447_), .A3(new_n434_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n449_), .B1(new_n462_), .B2(new_n423_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n395_), .B(new_n459_), .C1(new_n463_), .C2(new_n435_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n420_), .A2(new_n421_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n422_), .B1(new_n460_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n459_), .B1(new_n463_), .B2(new_n435_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n405_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n422_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n465_), .A4(new_n464_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(KEYINPUT73), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G190gat), .B(G218gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT72), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G134gat), .B(G162gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(KEYINPUT36), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n467_), .A2(KEYINPUT73), .A3(new_n471_), .A4(new_n477_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(KEYINPUT36), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT74), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT37), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G231gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT77), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n392_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G57gat), .B(G64gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT11), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT68), .B(G71gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(new_n284_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n493_), .B(G78gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n490_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G127gat), .B(G155gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT16), .ZN(new_n503_));
  XOR2_X1   g302(.A(G183gat), .B(G211gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n490_), .A2(new_n500_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n501_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n505_), .B(KEYINPUT17), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n483_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n486_), .A2(KEYINPUT37), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n486_), .A2(KEYINPUT37), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n499_), .B(new_n459_), .C1(new_n463_), .C2(new_n435_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n468_), .A2(new_n500_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n468_), .B2(new_n500_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n520_), .B(new_n521_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n468_), .A2(new_n500_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n518_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n521_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n525_), .A2(new_n529_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(KEYINPUT70), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(new_n537_), .A3(new_n540_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n525_), .A2(new_n529_), .A3(new_n536_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n536_), .B1(new_n525_), .B2(new_n529_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n487_), .A2(new_n513_), .A3(new_n517_), .A4(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n383_), .A2(new_n417_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n384_), .A3(new_n362_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT38), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT99), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n380_), .A2(new_n381_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n362_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n378_), .A3(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n371_), .A2(new_n360_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n300_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n514_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT100), .ZN(new_n560_));
  INV_X1    g359(.A(new_n546_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(new_n417_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n513_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n559_), .B2(KEYINPUT100), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(G1gat), .B1(new_n565_), .B2(new_n555_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n552_), .A2(new_n553_), .A3(new_n566_), .ZN(G1324gat));
  NAND3_X1  g366(.A1(new_n548_), .A2(new_n385_), .A3(new_n377_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n560_), .A2(new_n564_), .A3(new_n377_), .A4(new_n562_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT39), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(G8gat), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n569_), .B2(G8gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n568_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(KEYINPUT40), .B(new_n568_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(G1325gat));
  OAI21_X1  g377(.A(G15gat), .B1(new_n565_), .B2(new_n248_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT41), .Z(new_n580_));
  INV_X1    g379(.A(G15gat), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n548_), .A2(new_n581_), .A3(new_n247_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(G1326gat));
  INV_X1    g382(.A(G22gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n299_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n548_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G22gat), .B1(new_n565_), .B2(new_n299_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT42), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n587_), .A2(KEYINPUT42), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n586_), .B1(new_n589_), .B2(new_n590_), .ZN(G1327gat));
  NOR3_X1   g390(.A1(new_n561_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n558_), .A2(new_n416_), .A3(new_n592_), .ZN(new_n593_));
  OR3_X1    g392(.A1(new_n593_), .A2(G29gat), .A3(new_n555_), .ZN(new_n594_));
  AND4_X1   g393(.A1(new_n515_), .A2(new_n481_), .A3(new_n484_), .A4(new_n516_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n516_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n558_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT43), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n513_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n558_), .A2(KEYINPUT43), .A3(new_n598_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n562_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT44), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n601_), .A2(KEYINPUT44), .A3(new_n562_), .A4(new_n602_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n362_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G29gat), .B1(new_n607_), .B2(new_n608_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n594_), .B1(new_n609_), .B2(new_n610_), .ZN(G1328gat));
  NAND3_X1  g410(.A1(new_n605_), .A2(new_n377_), .A3(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G36gat), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n593_), .A2(G36gat), .A3(new_n378_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT45), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT46), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(new_n615_), .A3(KEYINPUT46), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1329gat));
  NAND4_X1  g419(.A1(new_n605_), .A2(G43gat), .A3(new_n247_), .A4(new_n606_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT102), .B(G43gat), .Z(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n593_), .B2(new_n248_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g424(.A1(new_n593_), .A2(new_n299_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(G50gat), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n605_), .A2(new_n606_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n585_), .A2(G50gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(G1331gat));
  AND2_X1   g429(.A1(new_n560_), .A2(new_n564_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n546_), .A2(new_n416_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n362_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G57gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n383_), .A2(new_n416_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n597_), .A2(new_n513_), .A3(new_n561_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n636_), .A2(KEYINPUT103), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(KEYINPUT103), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n555_), .A2(G57gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n634_), .B1(new_n639_), .B2(new_n640_), .ZN(G1332gat));
  OR3_X1    g440(.A1(new_n639_), .A2(G64gat), .A3(new_n378_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n631_), .A2(new_n377_), .A3(new_n632_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(G64gat), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n643_), .B2(G64gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(G1333gat));
  OR3_X1    g447(.A1(new_n639_), .A2(G71gat), .A3(new_n248_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n631_), .A2(new_n247_), .A3(new_n632_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT49), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(G71gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n650_), .B2(G71gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n649_), .B1(new_n653_), .B2(new_n654_), .ZN(G1334gat));
  NAND3_X1  g454(.A1(new_n631_), .A2(new_n585_), .A3(new_n632_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(G78gat), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n656_), .B2(G78gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n585_), .A2(new_n284_), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n659_), .A2(new_n660_), .B1(new_n639_), .B2(new_n661_), .ZN(G1335gat));
  NOR3_X1   g461(.A1(new_n513_), .A2(new_n546_), .A3(new_n514_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n635_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G85gat), .B1(new_n664_), .B2(new_n362_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT106), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n601_), .A2(new_n602_), .A3(new_n632_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n667_), .A2(new_n555_), .A3(new_n452_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1336gat));
  OAI21_X1  g468(.A(G92gat), .B1(new_n667_), .B2(new_n378_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n664_), .A2(new_n453_), .A3(new_n377_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1337gat));
  NAND4_X1  g471(.A1(new_n601_), .A2(new_n247_), .A3(new_n602_), .A4(new_n632_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n247_), .A2(new_n456_), .ZN(new_n674_));
  AOI22_X1  g473(.A1(new_n673_), .A2(G99gat), .B1(new_n664_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(KEYINPUT51), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(KEYINPUT51), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n678_), .B(new_n679_), .Z(G1338gat));
  NAND3_X1  g479(.A1(new_n664_), .A2(new_n457_), .A3(new_n585_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n601_), .A2(new_n585_), .A3(new_n602_), .A4(new_n632_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT52), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G106gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G106gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g486(.A(KEYINPUT54), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n547_), .A2(new_n416_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n693_));
  NOR4_X1   g492(.A1(new_n547_), .A2(KEYINPUT108), .A3(KEYINPUT109), .A4(new_n416_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n597_), .A2(new_n417_), .A3(new_n513_), .A4(new_n546_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT109), .B1(new_n696_), .B2(KEYINPUT108), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT54), .B1(new_n696_), .B2(KEYINPUT108), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n689_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n695_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT56), .ZN(new_n702_));
  INV_X1    g501(.A(new_n522_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n526_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n468_), .A2(new_n500_), .A3(new_n522_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n706_), .A2(KEYINPUT55), .A3(new_n521_), .A4(new_n520_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n520_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n528_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT55), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n525_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n525_), .A2(KEYINPUT110), .A3(new_n711_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n702_), .B1(new_n716_), .B2(new_n536_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n536_), .A2(new_n702_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT111), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n715_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT110), .B1(new_n525_), .B2(new_n711_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n707_), .B(new_n709_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n718_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n717_), .A2(new_n720_), .A3(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n417_), .A2(new_n542_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n399_), .A2(new_n400_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n412_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n401_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT112), .B1(new_n732_), .B2(new_n414_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n397_), .A2(new_n406_), .A3(new_n401_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n415_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n544_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n485_), .B1(new_n728_), .B2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n415_), .A3(new_n537_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n723_), .A2(new_n718_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n717_), .B2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT58), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n597_), .B1(new_n742_), .B2(KEYINPUT58), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n739_), .A2(KEYINPUT57), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n737_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n485_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n746_), .C1(new_n747_), .C2(new_n485_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n749_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n701_), .B1(new_n752_), .B2(new_n563_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n555_), .A2(new_n377_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n299_), .A3(new_n247_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(new_n755_), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT114), .B1(new_n753_), .B2(new_n757_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(G113gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n416_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT59), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n757_), .B2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n765_), .B2(new_n757_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n747_), .A2(new_n746_), .A3(new_n485_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n743_), .A2(new_n744_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n748_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n748_), .A2(new_n769_), .A3(KEYINPUT116), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n513_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n767_), .B1(new_n774_), .B2(new_n701_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT59), .B1(new_n753_), .B2(new_n757_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT117), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT117), .B1(new_n775_), .B2(new_n776_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n417_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n763_), .B1(new_n779_), .B2(new_n762_), .ZN(G1340gat));
  NAND3_X1  g579(.A1(new_n775_), .A2(new_n776_), .A3(new_n561_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT118), .B(G120gat), .Z(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n782_), .A2(KEYINPUT60), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n546_), .B2(KEYINPUT60), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n759_), .A2(new_n760_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n784_), .A2(new_n790_), .A3(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1341gat));
  AOI21_X1  g591(.A(G127gat), .B1(new_n761_), .B2(new_n513_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n777_), .A2(new_n778_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n513_), .A2(G127gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT120), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n794_), .B2(new_n796_), .ZN(G1342gat));
  INV_X1    g596(.A(G134gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n761_), .A2(new_n798_), .A3(new_n485_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n777_), .A2(new_n778_), .A3(new_n597_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n798_), .ZN(G1343gat));
  NOR4_X1   g600(.A1(new_n753_), .A2(new_n377_), .A3(new_n555_), .A4(new_n380_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n416_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n561_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n513_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT61), .B(G155gat), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(G1346gat));
  INV_X1    g608(.A(G162gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n802_), .A2(new_n810_), .A3(new_n485_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n802_), .A2(new_n598_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n810_), .ZN(G1347gat));
  NOR2_X1   g612(.A1(new_n774_), .A2(new_n701_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n555_), .A2(new_n377_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n248_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n416_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT121), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n299_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G169gat), .B1(new_n814_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT62), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n814_), .A2(new_n381_), .A3(new_n815_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n416_), .A3(new_n305_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1348gat));
  NAND3_X1  g623(.A1(new_n816_), .A2(G176gat), .A3(new_n561_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n753_), .A2(new_n585_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n561_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n211_), .ZN(G1349gat));
  AND2_X1   g627(.A1(new_n513_), .A2(new_n302_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n754_), .A2(new_n299_), .A3(new_n513_), .A4(new_n816_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n822_), .A2(new_n829_), .B1(new_n208_), .B2(new_n830_), .ZN(G1350gat));
  NAND2_X1  g630(.A1(new_n822_), .A2(new_n598_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G190gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n822_), .A2(new_n225_), .A3(new_n485_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1351gat));
  NOR2_X1   g634(.A1(new_n380_), .A2(new_n362_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(KEYINPUT122), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(KEYINPUT122), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n378_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n754_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n416_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n546_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G204gat), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT123), .B(G204gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n844_), .B2(new_n848_), .ZN(G1353gat));
  OAI22_X1  g648(.A1(new_n840_), .A2(new_n563_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT63), .B(G211gat), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n754_), .A2(new_n839_), .A3(new_n513_), .A4(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1354gat));
  INV_X1    g656(.A(KEYINPUT126), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT125), .B(G218gat), .Z(new_n859_));
  AND3_X1   g658(.A1(new_n841_), .A2(new_n598_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n841_), .B2(new_n485_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n841_), .A2(new_n598_), .A3(new_n859_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n840_), .A2(new_n514_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n863_), .B(KEYINPUT126), .C1(new_n864_), .C2(new_n859_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1355gat));
endmodule


