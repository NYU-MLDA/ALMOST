//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  OR3_X1    g003(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT66), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(KEYINPUT66), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT8), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G92gat), .Z(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n212_), .A2(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT10), .B(G99gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(new_n203_), .C1(G106gat), .C2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n210_), .A2(KEYINPUT8), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n211_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G71gat), .B(G78gat), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(new_n226_), .A3(KEYINPUT11), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT12), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G230gat), .A2(G233gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n211_), .A2(new_n221_), .A3(new_n229_), .A4(new_n220_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n222_), .A2(KEYINPUT12), .A3(new_n230_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n235_), .B(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n230_), .B2(new_n222_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n237_), .B1(new_n240_), .B2(new_n234_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G120gat), .B(G148gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT69), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G176gat), .B(G204gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n237_), .B(new_n247_), .C1(new_n240_), .C2(new_n234_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT13), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n249_), .A2(new_n250_), .B1(KEYINPUT70), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT37), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G232gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT34), .Z(new_n259_));
  XNOR2_X1  g058(.A(G29gat), .B(G36gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G43gat), .B(G50gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n222_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n262_), .B(KEYINPUT15), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n222_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n259_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G162gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT73), .B(G134gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT36), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n282_), .B(KEYINPUT74), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(KEYINPUT75), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n277_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n281_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(KEYINPUT36), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n275_), .A2(new_n276_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n257_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI211_X1 g096(.A(KEYINPUT76), .B(new_n257_), .C1(new_n291_), .C2(new_n294_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n294_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n284_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT37), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n297_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT102), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT87), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n308_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n308_), .A3(KEYINPUT87), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT2), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321_));
  INV_X1    g120(.A(G141gat), .ZN(new_n322_));
  INV_X1    g121(.A(G148gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n315_), .B1(new_n320_), .B2(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n317_), .A2(new_n319_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n331_), .A2(KEYINPUT88), .A3(new_n325_), .A4(new_n324_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT89), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n328_), .A2(KEYINPUT1), .B1(new_n322_), .B2(new_n323_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n316_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n333_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n334_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n314_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n309_), .A2(new_n311_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n342_), .A3(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT97), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT97), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n333_), .A2(new_n345_), .A3(new_n342_), .A4(new_n338_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n306_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n314_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n333_), .A2(new_n338_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT89), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n333_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n349_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT4), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n305_), .B1(new_n348_), .B2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n344_), .A2(new_n346_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n356_), .A2(new_n353_), .A3(new_n305_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(new_n212_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT0), .B(G57gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n355_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT101), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n355_), .A2(new_n358_), .A3(new_n366_), .A4(new_n363_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n303_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT28), .B(G22gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n351_), .A2(new_n352_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n373_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n374_));
  INV_X1    g173(.A(G50gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n339_), .A2(new_n340_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n372_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(G50gat), .B1(new_n373_), .B2(KEYINPUT29), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n377_), .A3(new_n375_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n371_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT93), .ZN(new_n384_));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387_));
  INV_X1    g186(.A(G197gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G204gat), .ZN(new_n389_));
  INV_X1    g188(.A(G204gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G197gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(KEYINPUT21), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n390_), .B2(G197gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n391_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(KEYINPUT21), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n398_), .B2(KEYINPUT21), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n387_), .B(new_n394_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n387_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(KEYINPUT21), .A3(new_n392_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n408_));
  AOI211_X1 g207(.A(KEYINPUT92), .B(new_n377_), .C1(new_n333_), .C2(new_n338_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n403_), .A2(new_n405_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n411_), .B(new_n413_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n386_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n384_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n414_), .B(new_n385_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n383_), .A3(KEYINPUT93), .A4(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n383_), .A2(new_n419_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT4), .B1(new_n356_), .B2(new_n353_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n341_), .A2(new_n306_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n304_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n362_), .B1(new_n426_), .B2(new_n357_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n355_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(KEYINPUT101), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(KEYINPUT102), .A3(new_n368_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n370_), .A2(new_n423_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT100), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT25), .B(G183gat), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT83), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT25), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT83), .B1(new_n435_), .B2(G183gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT84), .B(G190gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT26), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n434_), .B(new_n436_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G169gat), .ZN(new_n442_));
  INV_X1    g241(.A(G176gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT85), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(G169gat), .B2(G176gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n444_), .A2(new_n446_), .A3(KEYINPUT24), .A4(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G183gat), .A2(G190gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT23), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT24), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n445_), .A2(G169gat), .A3(G176gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT85), .B1(new_n442_), .B2(new_n443_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n441_), .A2(new_n451_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G183gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n437_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n450_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n447_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT22), .B(G169gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n443_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n456_), .A2(new_n403_), .A3(new_n463_), .A4(new_n405_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT26), .B(G190gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n433_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n451_), .A2(KEYINPUT95), .A3(new_n455_), .A4(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n455_), .A2(new_n466_), .A3(new_n450_), .A4(new_n448_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT95), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n450_), .B1(G183gat), .B2(G190gat), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n467_), .A2(new_n470_), .B1(new_n462_), .B2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n464_), .B(KEYINPUT20), .C1(new_n406_), .C2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n432_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n462_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n468_), .A2(new_n469_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n468_), .A2(new_n469_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n479_), .B1(new_n483_), .B2(new_n413_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n484_), .A2(KEYINPUT100), .A3(new_n476_), .A4(new_n464_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n406_), .A2(new_n480_), .A3(new_n468_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n456_), .A2(new_n463_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n479_), .B1(new_n487_), .B2(new_n413_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n478_), .B(new_n485_), .C1(new_n476_), .C2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G8gat), .B(G36gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G92gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT18), .B(G64gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n477_), .B1(new_n406_), .B2(new_n472_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n473_), .A2(new_n477_), .B1(new_n497_), .B2(new_n488_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n494_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(KEYINPUT27), .A3(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT96), .B1(new_n498_), .B2(new_n494_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT96), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n497_), .A2(new_n488_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n476_), .B1(new_n484_), .B2(new_n464_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n502_), .B(new_n495_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n505_), .A3(new_n499_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT103), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT27), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n500_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT104), .B1(new_n431_), .B2(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n429_), .A2(KEYINPUT102), .A3(new_n368_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT102), .B1(new_n429_), .B2(new_n368_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT104), .ZN(new_n517_));
  INV_X1    g316(.A(new_n500_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n506_), .A2(new_n508_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT103), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n520_), .B2(new_n509_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n516_), .A2(new_n517_), .A3(new_n423_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n498_), .ZN(new_n523_));
  OAI211_X1 g322(.A(KEYINPUT32), .B(new_n494_), .C1(new_n523_), .C2(KEYINPUT99), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(new_n490_), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n498_), .A2(KEYINPUT99), .B1(KEYINPUT32), .B2(new_n494_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n368_), .B(new_n429_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n364_), .B(KEYINPUT33), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n341_), .A2(new_n347_), .A3(new_n305_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n529_), .A2(new_n362_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT98), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n304_), .B1(new_n348_), .B2(new_n354_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(KEYINPUT98), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n534_), .A2(new_n499_), .A3(new_n501_), .A4(new_n505_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n527_), .B1(new_n528_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n422_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n513_), .A2(new_n522_), .A3(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n314_), .B(KEYINPUT30), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n487_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G15gat), .B(G43gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G71gat), .B(G99gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n540_), .A2(new_n543_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n538_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n551_), .A2(new_n422_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT105), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT105), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n554_), .A2(new_n516_), .A3(new_n557_), .A4(new_n521_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(G1gat), .ZN(new_n564_));
  INV_X1    g363(.A(G8gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT77), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G15gat), .B(G22gat), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT77), .B(KEYINPUT14), .C1(new_n564_), .C2(new_n565_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G1gat), .B(G8gat), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n572_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n263_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(new_n574_), .A3(new_n262_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(G229gat), .A3(G233gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n269_), .A2(new_n575_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n577_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n579_), .A2(KEYINPUT80), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT80), .B1(new_n579_), .B2(new_n582_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n563_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT81), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n579_), .A2(new_n582_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n563_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n586_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n588_), .A2(new_n592_), .A3(KEYINPUT82), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT82), .B1(new_n588_), .B2(new_n592_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n560_), .A2(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT106), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT106), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n256_), .B(new_n302_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n575_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n230_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n602_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT79), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n602_), .A2(new_n608_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(KEYINPUT17), .B2(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n599_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n516_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n564_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n538_), .A2(new_n552_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n299_), .A2(new_n300_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n613_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n595_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n256_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n516_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n616_), .A2(KEYINPUT38), .A3(new_n564_), .A4(new_n617_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(new_n627_), .A3(new_n628_), .ZN(G1324gat));
  NAND2_X1  g428(.A1(new_n512_), .A2(new_n565_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G8gat), .B1(new_n626_), .B2(new_n521_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(KEYINPUT39), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(KEYINPUT39), .ZN(new_n633_));
  OAI22_X1  g432(.A1(new_n615_), .A2(new_n630_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n626_), .B2(new_n552_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT41), .Z(new_n638_));
  OR2_X1    g437(.A1(new_n615_), .A2(G15gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n552_), .ZN(G1326gat));
  OAI21_X1  g439(.A(G22gat), .B1(new_n626_), .B2(new_n422_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT42), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n615_), .A2(G22gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(new_n422_), .ZN(G1327gat));
  NAND2_X1  g443(.A1(new_n597_), .A2(new_n598_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n256_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n622_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n614_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n617_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n560_), .B2(new_n302_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n286_), .B(new_n289_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT37), .B1(new_n653_), .B2(new_n299_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT76), .ZN(new_n655_));
  INV_X1    g454(.A(new_n301_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n295_), .A2(new_n296_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n621_), .A2(KEYINPUT43), .A3(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n625_), .B(new_n613_), .C1(new_n652_), .C2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n560_), .A2(new_n651_), .A3(new_n302_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n621_), .B2(new_n658_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n625_), .A4(new_n613_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n617_), .A2(G29gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n650_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n649_), .A2(KEYINPUT45), .A3(new_n670_), .A4(new_n512_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n662_), .A2(new_n512_), .A3(new_n666_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G36gat), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n645_), .A2(new_n670_), .A3(new_n646_), .A4(new_n648_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(new_n521_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n671_), .A2(new_n673_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n671_), .A2(KEYINPUT46), .A3(new_n676_), .A4(new_n673_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  AND2_X1   g480(.A1(new_n551_), .A2(G43gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n662_), .A2(new_n666_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n662_), .A2(KEYINPUT107), .A3(new_n666_), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT108), .B(G43gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n552_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT47), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n687_), .A2(new_n693_), .A3(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1330gat));
  AOI21_X1  g494(.A(G50gat), .B1(new_n649_), .B2(new_n423_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n422_), .A2(new_n375_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n667_), .B2(new_n697_), .ZN(G1331gat));
  NAND3_X1  g497(.A1(new_n658_), .A2(new_n256_), .A3(new_n614_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT109), .Z(new_n700_));
  NOR2_X1   g499(.A1(new_n621_), .A2(new_n595_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n617_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT110), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n623_), .A2(new_n624_), .A3(new_n256_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT111), .B(G57gat), .Z(new_n706_));
  NOR3_X1   g505(.A1(new_n705_), .A2(new_n516_), .A3(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1332gat));
  OAI21_X1  g507(.A(G64gat), .B1(new_n705_), .B2(new_n521_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  INV_X1    g509(.A(new_n702_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n521_), .A2(G64gat), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT112), .Z(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n711_), .B2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n705_), .B2(new_n552_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n711_), .A2(G71gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n552_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n705_), .B2(new_n422_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n711_), .A2(G78gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n422_), .ZN(G1335gat));
  NAND2_X1  g521(.A1(new_n256_), .A2(new_n624_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n621_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n648_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n617_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n723_), .A2(new_n614_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n665_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT113), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n665_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n516_), .A2(new_n212_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n727_), .B1(new_n733_), .B2(new_n734_), .ZN(G1336gat));
  AOI21_X1  g534(.A(G92gat), .B1(new_n726_), .B2(new_n512_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n521_), .A2(new_n213_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n733_), .B2(new_n737_), .ZN(G1337gat));
  NOR3_X1   g537(.A1(new_n725_), .A2(new_n219_), .A3(new_n552_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n730_), .A2(new_n551_), .A3(new_n732_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G99gat), .ZN(new_n741_));
  OR2_X1    g540(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n742_));
  NAND2_X1  g541(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1338gat));
  OAI211_X1 g545(.A(new_n423_), .B(new_n728_), .C1(new_n652_), .C2(new_n659_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT115), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n665_), .A2(new_n749_), .A3(new_n423_), .A4(new_n728_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(G106gat), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT52), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n748_), .A2(new_n753_), .A3(G106gat), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n725_), .A2(G106gat), .A3(new_n422_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  NOR2_X1   g560(.A1(new_n516_), .A2(new_n512_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n554_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n234_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n233_), .A2(new_n236_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n239_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n222_), .A2(KEYINPUT12), .A3(new_n230_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT12), .B1(new_n222_), .B2(new_n230_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT55), .A3(new_n234_), .A4(new_n235_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n237_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n766_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n248_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT117), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n595_), .A3(new_n250_), .A4(new_n778_), .ZN(new_n779_));
  AND4_X1   g578(.A1(G229gat), .A2(new_n580_), .A3(G233gat), .A4(new_n577_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n581_), .B2(new_n578_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n590_), .B1(new_n781_), .B2(new_n563_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n251_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n779_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n647_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n774_), .A2(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n773_), .A2(new_n776_), .A3(new_n248_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n250_), .A2(new_n782_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT118), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n250_), .A2(new_n782_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n790_), .A2(KEYINPUT58), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n795_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n790_), .A2(new_n795_), .A3(KEYINPUT119), .A4(KEYINPUT58), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n302_), .A2(new_n798_), .A3(new_n801_), .A4(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n784_), .A2(KEYINPUT57), .A3(new_n647_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n787_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n784_), .B2(new_n647_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n786_), .B(new_n622_), .C1(new_n779_), .C2(new_n783_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT120), .A3(new_n803_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n811_), .A3(new_n613_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n595_), .B2(new_n613_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n624_), .A2(KEYINPUT116), .A3(new_n614_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n658_), .A2(new_n646_), .A3(new_n814_), .A4(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT54), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n763_), .B1(new_n812_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n595_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n812_), .A2(new_n817_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n763_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT59), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n805_), .A2(new_n613_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n817_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n821_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n595_), .A2(G113gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n819_), .B1(new_n828_), .B2(new_n829_), .ZN(G1340gat));
  NAND4_X1  g629(.A1(new_n823_), .A2(KEYINPUT121), .A3(new_n256_), .A4(new_n827_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n256_), .B(new_n827_), .C1(new_n818_), .C2(new_n826_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(G120gat), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n646_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n818_), .B(new_n837_), .C1(KEYINPUT60), .C2(new_n836_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(G1341gat));
  AOI21_X1  g638(.A(G127gat), .B1(new_n818_), .B2(new_n614_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n614_), .A2(G127gat), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n828_), .B2(new_n842_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n822_), .B2(new_n647_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n658_), .A2(new_n844_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n827_), .B(new_n846_), .C1(new_n818_), .C2(new_n826_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT122), .ZN(G1343gat));
  AOI211_X1 g648(.A(new_n551_), .B(new_n422_), .C1(new_n812_), .C2(new_n817_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n762_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n624_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT123), .B(G141gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n851_), .A2(new_n646_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n323_), .ZN(G1345gat));
  NOR2_X1   g655(.A1(new_n851_), .A2(new_n613_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT61), .B(G155gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n851_), .A2(new_n860_), .A3(new_n658_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n850_), .A2(new_n622_), .A3(new_n762_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(new_n862_), .ZN(G1347gat));
  NOR2_X1   g662(.A1(new_n617_), .A2(new_n521_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n554_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n614_), .B1(new_n810_), .B2(new_n803_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n816_), .B(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n595_), .B(new_n866_), .C1(new_n867_), .C2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n825_), .A2(KEYINPUT124), .A3(new_n595_), .A4(new_n866_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(G169gat), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n825_), .A2(new_n866_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n595_), .A3(new_n461_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n872_), .A2(new_n873_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n876_), .A2(KEYINPUT125), .A3(new_n879_), .A4(new_n880_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1348gat));
  AOI21_X1  g684(.A(G176gat), .B1(new_n878_), .B2(new_n256_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n865_), .B1(new_n812_), .B2(new_n817_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n646_), .A2(new_n443_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  AOI21_X1  g688(.A(G183gat), .B1(new_n887_), .B2(new_n614_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n613_), .A2(new_n433_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n878_), .B2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n877_), .B2(new_n658_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n622_), .A2(new_n465_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT126), .Z(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n877_), .B2(new_n896_), .ZN(G1351gat));
  NAND2_X1  g696(.A1(new_n850_), .A2(new_n864_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n624_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n388_), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n646_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT127), .B(G204gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1353gat));
  INV_X1    g702(.A(new_n898_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT63), .B(G211gat), .Z(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n614_), .A3(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n898_), .B2(new_n613_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1354gat));
  AND3_X1   g708(.A1(new_n904_), .A2(G218gat), .A3(new_n302_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G218gat), .B1(new_n904_), .B2(new_n622_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1355gat));
endmodule


