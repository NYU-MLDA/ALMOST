//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n971_,
    new_n972_, new_n973_, new_n975_, new_n976_, new_n978_, new_n979_,
    new_n980_, new_n982_, new_n983_, new_n984_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_,
    new_n995_;
  INV_X1    g000(.A(G50gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G29gat), .A2(G36gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT69), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n206_));
  AND2_X1   g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G43gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n205_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n205_), .B2(new_n209_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n202_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n207_), .A2(new_n208_), .A3(new_n206_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT69), .B1(new_n203_), .B2(new_n204_), .ZN(new_n215_));
  OAI21_X1  g014(.A(G43gat), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n205_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(G50gat), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n213_), .A2(new_n218_), .A3(KEYINPUT15), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT6), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT6), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n224_), .B(new_n228_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G85gat), .B(G92gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT8), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n238_), .A3(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(KEYINPUT9), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT10), .B(G99gat), .Z(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n227_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n231_), .A2(KEYINPUT6), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n229_), .A2(G99gat), .A3(G106gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G85gat), .ZN(new_n247_));
  INV_X1    g046(.A(G92gat), .ZN(new_n248_));
  OR3_X1    g047(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT9), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n241_), .A2(new_n243_), .A3(new_n246_), .A4(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT65), .B1(new_n240_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n224_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI211_X1 g053(.A(KEYINPUT8), .B(new_n234_), .C1(new_n254_), .C2(new_n246_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n238_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n256_));
  OAI211_X1 g055(.A(KEYINPUT65), .B(new_n250_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n223_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n250_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(new_n219_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT34), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(KEYINPUT35), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(KEYINPUT35), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n264_), .A2(KEYINPUT35), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n259_), .A2(new_n266_), .A3(new_n267_), .A4(new_n261_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G134gat), .ZN(new_n271_));
  INV_X1    g070(.A(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT36), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT37), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n273_), .B(KEYINPUT36), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT70), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n276_), .A2(new_n277_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n269_), .A2(new_n278_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n276_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n269_), .A2(KEYINPUT71), .A3(new_n278_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n287_), .B2(new_n277_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G71gat), .B(G78gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(G57gat), .B(G64gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT11), .A3(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(G57gat), .A2(G64gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G57gat), .A2(G64gat), .ZN(new_n294_));
  OR3_X1    g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT11), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT11), .B1(new_n293_), .B2(new_n294_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G71gat), .B(G78gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n292_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT72), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G8gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n305_), .A3(G1gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT14), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT73), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n309_), .A3(KEYINPUT14), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n302_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n306_), .A2(new_n309_), .A3(KEYINPUT14), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n309_), .B1(new_n306_), .B2(KEYINPUT14), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n302_), .B(new_n312_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n301_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n312_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G1gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G8gat), .A3(new_n316_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G231gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n322_), .A2(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n300_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n299_), .A3(new_n325_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT75), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G127gat), .B(G155gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G183gat), .B(G211gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n331_), .A2(KEYINPUT17), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n328_), .A2(new_n330_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n337_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(KEYINPUT17), .C1(new_n331_), .C2(new_n337_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n289_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT76), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT84), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT87), .ZN(new_n349_));
  INV_X1    g148(.A(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(G169gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n351_), .A2(KEYINPUT22), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n350_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n347_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT88), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT23), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n357_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT79), .B(G183gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(G190gat), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n363_), .B(new_n347_), .C1(new_n349_), .C2(new_n354_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n356_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n351_), .A2(new_n350_), .A3(KEYINPUT83), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(G169gat), .B2(G176gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n347_), .A3(KEYINPUT24), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT85), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n370_), .A2(new_n347_), .A3(new_n373_), .A4(KEYINPUT24), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n357_), .A2(KEYINPUT23), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n359_), .B2(new_n357_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n361_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n361_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT26), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(KEYINPUT82), .B2(G190gat), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n382_), .A2(KEYINPUT81), .ZN(new_n386_));
  INV_X1    g185(.A(G183gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(KEYINPUT81), .B2(new_n382_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(KEYINPUT82), .A3(G190gat), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n380_), .A2(new_n383_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n369_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n365_), .B1(new_n378_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G197gat), .B(G204gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT95), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT21), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n396_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n402_), .A2(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n397_), .A2(KEYINPUT21), .A3(new_n398_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n401_), .A2(KEYINPUT96), .A3(new_n403_), .A4(new_n404_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n395_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT19), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n345_), .A2(KEYINPUT24), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n414_), .A2(KEYINPUT100), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(KEYINPUT100), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n370_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT25), .B(G183gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n384_), .A2(G190gat), .ZN(new_n419_));
  INV_X1    g218(.A(G190gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT26), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n419_), .A2(new_n421_), .A3(KEYINPUT99), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT99), .B1(new_n419_), .B2(new_n421_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n418_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n417_), .A2(new_n424_), .A3(new_n393_), .A4(new_n360_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n348_), .A2(new_n350_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G183gat), .A2(G190gat), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n347_), .B(new_n426_), .C1(new_n376_), .C2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n405_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n410_), .A2(KEYINPUT20), .A3(new_n413_), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n428_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n404_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT21), .B1(new_n397_), .B2(new_n398_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n403_), .A3(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT20), .B(new_n435_), .C1(new_n395_), .C2(new_n409_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n436_), .A2(KEYINPUT101), .A3(new_n412_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT101), .B1(new_n436_), .B2(new_n412_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n430_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT18), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G64gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(new_n248_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n443_), .B(new_n430_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT27), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n436_), .A2(new_n412_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n449_), .A2(KEYINPUT102), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(KEYINPUT102), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n429_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n413_), .B1(new_n410_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n444_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(KEYINPUT27), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G120gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G127gat), .B(G134gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT89), .ZN(new_n459_));
  INV_X1    g258(.A(G113gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(G127gat), .A2(G134gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G127gat), .A2(G134gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n459_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n460_), .B1(new_n459_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n457_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n459_), .A2(new_n464_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G113gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n459_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(G120gat), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT1), .ZN(new_n474_));
  INV_X1    g273(.A(G155gat), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n474_), .A2(KEYINPUT91), .B1(new_n475_), .B2(new_n272_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n477_), .A3(KEYINPUT1), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n473_), .B2(KEYINPUT1), .ZN(new_n480_));
  OR3_X1    g279(.A1(new_n473_), .A2(new_n479_), .A3(KEYINPUT1), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n476_), .A2(new_n478_), .A3(new_n480_), .A4(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G141gat), .A2(G148gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT90), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G141gat), .A2(G148gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n475_), .A2(new_n272_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n473_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT2), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n483_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n485_), .B(KEYINPUT3), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n489_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT93), .B1(new_n487_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n491_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n483_), .B(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n493_), .B(new_n496_), .C1(new_n498_), .C2(KEYINPUT2), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n488_), .A3(new_n473_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n482_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT93), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n472_), .B1(new_n495_), .B2(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n472_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G29gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G85gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT0), .ZN(new_n512_));
  INV_X1    g311(.A(G57gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n504_), .A2(KEYINPUT4), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n495_), .A2(new_n503_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n472_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n472_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n515_), .B1(new_n520_), .B2(KEYINPUT4), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n509_), .B(new_n514_), .C1(new_n521_), .C2(new_n506_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n514_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT4), .B1(new_n504_), .B2(new_n505_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n506_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n523_), .B1(new_n527_), .B2(new_n508_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n447_), .A2(new_n456_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G71gat), .B(G99gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT30), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G227gat), .A2(G233gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n395_), .A2(new_n472_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n395_), .A2(new_n472_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G15gat), .B(G43gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT31), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n536_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n517_), .B(new_n365_), .C1(new_n394_), .C2(new_n378_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n395_), .A2(new_n472_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n535_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n539_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n541_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n534_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n495_), .A2(new_n551_), .A3(new_n503_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G22gat), .B(G50gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT28), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n552_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G78gat), .B(G106gat), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n516_), .A2(KEYINPUT29), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G228gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT94), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n551_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n564_));
  OAI211_X1 g363(.A(G228gat), .B(G233gat), .C1(new_n564_), .C2(new_n405_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n558_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n557_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n551_), .B1(new_n495_), .B2(new_n503_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n561_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT96), .B1(new_n434_), .B2(new_n403_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n408_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n565_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n558_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n558_), .B(new_n565_), .C1(new_n569_), .C2(new_n573_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT97), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n550_), .B1(new_n568_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n567_), .B1(new_n566_), .B2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n556_), .B1(new_n576_), .B2(KEYINPUT97), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT98), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n557_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n549_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n545_), .A2(new_n548_), .ZN(new_n588_));
  AOI211_X1 g387(.A(new_n585_), .B(new_n588_), .C1(new_n579_), .C2(new_n583_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n530_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n591_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n529_), .B(new_n592_), .C1(new_n439_), .C2(new_n591_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n524_), .A2(new_n526_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n508_), .B1(new_n595_), .B2(new_n507_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n596_), .B2(new_n514_), .ZN(new_n597_));
  NOR4_X1   g396(.A1(new_n527_), .A2(new_n508_), .A3(KEYINPUT33), .A4(new_n523_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n446_), .B(new_n445_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n521_), .A2(new_n507_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n520_), .A2(new_n506_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n600_), .A2(new_n514_), .A3(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n593_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n568_), .A2(new_n578_), .A3(new_n550_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT98), .B1(new_n581_), .B2(new_n582_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n586_), .B(new_n588_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n590_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n219_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n321_), .ZN(new_n611_));
  AOI21_X1  g410(.A(G8gat), .B1(new_n320_), .B2(new_n316_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n223_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT78), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT78), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n613_), .A2(new_n614_), .A3(new_n618_), .A4(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT77), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n318_), .A2(new_n219_), .A3(new_n321_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n613_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n322_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(KEYINPUT77), .A3(new_n219_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n623_), .A2(new_n625_), .A3(G229gat), .A4(G233gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n620_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(new_n351_), .ZN(new_n629_));
  INV_X1    g428(.A(G197gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n631_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n620_), .A2(new_n626_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT13), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n299_), .B(new_n250_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT64), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT64), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n299_), .B1(new_n240_), .B2(new_n250_), .ZN(new_n640_));
  OR3_X1    g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT5), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(G176gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(G204gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT67), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n637_), .B1(new_n640_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n300_), .A2(KEYINPUT12), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT65), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n260_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(new_n257_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n651_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n649_), .B1(new_n656_), .B2(new_n642_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n652_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n650_), .B1(new_n260_), .B2(new_n300_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n637_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n659_), .A2(new_n662_), .A3(new_n649_), .A4(new_n642_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n644_), .B(new_n648_), .C1(new_n657_), .C2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT68), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n662_), .A3(new_n642_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT67), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n668_), .A2(new_n663_), .B1(new_n643_), .B2(new_n641_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT68), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n648_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n669_), .A2(new_n648_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n636_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n636_), .A3(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n609_), .A2(new_n635_), .A3(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n344_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n302_), .A3(new_n529_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT103), .Z(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT38), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT38), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n675_), .A2(new_n676_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n635_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT104), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n287_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n342_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n677_), .A2(new_n689_), .A3(new_n635_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n686_), .A2(new_n609_), .A3(new_n688_), .A4(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n529_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G1gat), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT105), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n682_), .A2(new_n683_), .A3(new_n694_), .ZN(G1324gat));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n447_), .A2(new_n456_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G8gat), .B1(new_n691_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT39), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n679_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n696_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n699_), .A2(new_n696_), .A3(new_n701_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT40), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n702_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1325gat));
  OAI21_X1  g508(.A(G15gat), .B1(new_n691_), .B2(new_n588_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT41), .Z(new_n711_));
  INV_X1    g510(.A(G15gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n679_), .A2(new_n712_), .A3(new_n549_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1326gat));
  OAI21_X1  g513(.A(new_n586_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT107), .Z(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G22gat), .B1(new_n691_), .B2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT42), .ZN(new_n719_));
  INV_X1    g518(.A(G22gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n679_), .A2(new_n720_), .A3(new_n716_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1327gat));
  NAND2_X1  g521(.A1(new_n342_), .A2(new_n687_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n678_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(G29gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n529_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n288_), .B1(new_n590_), .B2(new_n608_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT108), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT27), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n436_), .A2(new_n412_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n436_), .A2(KEYINPUT101), .A3(new_n412_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n443_), .B1(new_n735_), .B2(new_n430_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n446_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n730_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n692_), .A3(new_n455_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n715_), .A2(new_n588_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n584_), .A2(new_n586_), .A3(new_n549_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n736_), .A2(new_n737_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n602_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n743_), .B(new_n744_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n606_), .B1(new_n745_), .B2(new_n593_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n289_), .B1(new_n742_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(KEYINPUT43), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n727_), .A2(new_n728_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n729_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n686_), .A2(new_n342_), .A3(new_n690_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(KEYINPUT44), .A3(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n751_), .B2(new_n752_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n754_), .A2(new_n692_), .A3(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n726_), .B1(new_n756_), .B2(new_n725_), .ZN(G1328gat));
  NAND2_X1  g556(.A1(new_n751_), .A2(new_n752_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n697_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n753_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G36gat), .ZN(new_n763_));
  NOR4_X1   g562(.A1(new_n678_), .A2(G36gat), .A3(new_n697_), .A4(new_n723_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT45), .Z(new_n765_));
  OAI211_X1 g564(.A(new_n763_), .B(new_n765_), .C1(KEYINPUT109), .C2(KEYINPUT46), .ZN(new_n766_));
  NAND2_X1  g565(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1329gat));
  NAND3_X1  g567(.A1(new_n724_), .A2(new_n210_), .A3(new_n549_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n754_), .A2(new_n588_), .A3(new_n755_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n210_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g571(.A1(new_n760_), .A2(new_n715_), .A3(new_n753_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT110), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n760_), .A2(new_n775_), .A3(new_n715_), .A4(new_n753_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(G50gat), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n774_), .A2(KEYINPUT111), .A3(G50gat), .A4(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n716_), .A2(new_n202_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT112), .Z(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n724_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(G1331gat));
  INV_X1    g584(.A(new_n344_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n677_), .A2(new_n635_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n609_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(G57gat), .B1(new_n789_), .B2(new_n529_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n788_), .A2(new_n688_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n692_), .A2(new_n513_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n791_), .B2(new_n792_), .ZN(G1332gat));
  INV_X1    g592(.A(G64gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n791_), .B2(new_n761_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT48), .Z(new_n796_));
  NAND3_X1  g595(.A1(new_n789_), .A2(new_n794_), .A3(new_n761_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1333gat));
  INV_X1    g597(.A(G71gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n791_), .B2(new_n549_), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT49), .Z(new_n801_));
  NAND3_X1  g600(.A1(new_n789_), .A2(new_n799_), .A3(new_n549_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1334gat));
  INV_X1    g602(.A(G78gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n791_), .B2(new_n716_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT50), .Z(new_n806_));
  NAND3_X1  g605(.A1(new_n789_), .A2(new_n804_), .A3(new_n716_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1335gat));
  INV_X1    g607(.A(new_n723_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n788_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G85gat), .B1(new_n810_), .B2(new_n529_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n751_), .A2(new_n342_), .A3(new_n787_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n692_), .A2(new_n247_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(G1336gat));
  AOI21_X1  g613(.A(G92gat), .B1(new_n810_), .B2(new_n761_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n697_), .A2(new_n248_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n812_), .B2(new_n816_), .ZN(G1337gat));
  NAND3_X1  g616(.A1(new_n810_), .A2(new_n242_), .A3(new_n549_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT113), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n812_), .A2(new_n549_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G99gat), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT51), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(KEYINPUT51), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n824_), .B(new_n825_), .Z(G1338gat));
  NAND3_X1  g625(.A1(new_n810_), .A2(new_n227_), .A3(new_n715_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n751_), .A2(new_n715_), .A3(new_n342_), .A4(new_n787_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n828_), .A2(new_n829_), .A3(G106gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n828_), .B2(G106gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g632(.A1(new_n623_), .A2(new_n625_), .A3(new_n615_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n613_), .A2(new_n614_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n834_), .B(new_n631_), .C1(new_n835_), .C2(new_n615_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n634_), .A2(new_n836_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n837_), .A2(new_n672_), .A3(KEYINPUT116), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT116), .B1(new_n837_), .B2(new_n672_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT55), .B1(new_n668_), .B2(new_n663_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n667_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n656_), .A2(new_n642_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n840_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT56), .B1(new_n844_), .B2(new_n648_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n668_), .A2(new_n663_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n841_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n842_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n843_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  INV_X1    g650(.A(new_n648_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n845_), .A2(new_n853_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n838_), .A2(new_n839_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT58), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n837_), .A2(new_n672_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n844_), .A2(KEYINPUT56), .A3(new_n648_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n851_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n837_), .A2(new_n672_), .A3(KEYINPUT116), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(KEYINPUT117), .A3(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n857_), .A2(new_n289_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n843_), .B1(new_n846_), .B2(new_n841_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n648_), .B1(new_n869_), .B2(new_n848_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n851_), .B1(new_n870_), .B2(KEYINPUT115), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n632_), .A2(new_n634_), .B1(new_n666_), .B2(new_n671_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n873_), .B(KEYINPUT56), .C1(new_n844_), .C2(new_n648_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n872_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n672_), .A2(new_n673_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n837_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n878_), .B2(new_n287_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n880_), .B(new_n687_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n868_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n342_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n635_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n343_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n343_), .B2(new_n886_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n884_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n741_), .A2(new_n692_), .ZN(new_n892_));
  AND2_X1   g691(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n891_), .A2(new_n697_), .A3(new_n892_), .A4(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n342_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n868_), .B2(new_n882_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n697_), .B(new_n892_), .C1(new_n896_), .C2(new_n889_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n893_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n894_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n460_), .A2(KEYINPUT121), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n894_), .A2(new_n900_), .A3(KEYINPUT120), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT121), .B1(new_n685_), .B2(new_n460_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .A4(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n891_), .A2(new_n908_), .A3(new_n697_), .A4(new_n892_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n897_), .A2(KEYINPUT118), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n635_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n460_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n907_), .A2(new_n913_), .ZN(G1340gat));
  AOI21_X1  g713(.A(new_n457_), .B1(new_n901_), .B2(new_n684_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n457_), .A2(KEYINPUT60), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n457_), .B1(new_n677_), .B2(KEYINPUT60), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  AOI211_X1 g717(.A(new_n916_), .B(new_n918_), .C1(new_n909_), .C2(new_n910_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT122), .B1(new_n915_), .B2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n916_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n911_), .A2(new_n921_), .A3(new_n917_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n677_), .B1(new_n894_), .B2(new_n900_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n922_), .B(new_n923_), .C1(new_n457_), .C2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n920_), .A2(new_n925_), .ZN(G1341gat));
  AOI21_X1  g725(.A(G127gat), .B1(new_n911_), .B2(new_n895_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n903_), .A2(new_n905_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n895_), .A2(G127gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1342gat));
  AOI21_X1  g729(.A(G134gat), .B1(new_n911_), .B2(new_n687_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n289_), .A2(G134gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n928_), .B2(new_n932_), .ZN(G1343gat));
  NAND4_X1  g732(.A1(new_n891_), .A2(new_n529_), .A3(new_n587_), .A4(new_n697_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n635_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n684_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT123), .B1(new_n934_), .B2(new_n342_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n934_), .A2(KEYINPUT123), .A3(new_n342_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n941_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n944_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n946_), .A2(new_n940_), .A3(new_n942_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1346gat));
  NOR3_X1   g747(.A1(new_n934_), .A2(new_n272_), .A3(new_n288_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n935_), .A2(new_n687_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n272_), .B2(new_n950_), .ZN(G1347gat));
  NOR2_X1   g750(.A1(new_n697_), .A2(new_n529_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n549_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n717_), .B(new_n954_), .C1(new_n896_), .C2(new_n889_), .ZN(new_n955_));
  OAI21_X1  g754(.A(G169gat), .B1(new_n955_), .B2(new_n685_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n955_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n959_), .A2(new_n635_), .A3(new_n348_), .ZN(new_n960_));
  OAI211_X1 g759(.A(KEYINPUT62), .B(G169gat), .C1(new_n955_), .C2(new_n685_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n958_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(KEYINPUT124), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964_));
  NAND4_X1  g763(.A1(new_n958_), .A2(new_n960_), .A3(new_n964_), .A4(new_n961_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n965_), .ZN(G1348gat));
  AOI21_X1  g765(.A(G176gat), .B1(new_n959_), .B2(new_n684_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n891_), .A2(new_n586_), .A3(new_n584_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n968_), .A2(new_n350_), .A3(new_n677_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n967_), .B1(new_n969_), .B2(new_n954_), .ZN(G1349gat));
  NOR3_X1   g769(.A1(new_n955_), .A2(new_n418_), .A3(new_n342_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(KEYINPUT125), .ZN(new_n972_));
  OR3_X1    g771(.A1(new_n968_), .A2(new_n342_), .A3(new_n953_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n972_), .B1(new_n379_), .B2(new_n973_), .ZN(G1350gat));
  OAI21_X1  g773(.A(G190gat), .B1(new_n955_), .B2(new_n288_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n687_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n955_), .B2(new_n976_), .ZN(G1351gat));
  AOI21_X1  g776(.A(new_n740_), .B1(new_n884_), .B2(new_n890_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(new_n952_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n979_), .A2(new_n685_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(new_n980_), .B(new_n630_), .ZN(G1352gat));
  NOR2_X1   g780(.A1(new_n979_), .A2(new_n677_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n982_), .A2(KEYINPUT126), .A3(G204gat), .ZN(new_n983_));
  XOR2_X1   g782(.A(KEYINPUT126), .B(G204gat), .Z(new_n984_));
  AOI21_X1  g783(.A(new_n983_), .B1(new_n982_), .B2(new_n984_), .ZN(G1353gat));
  NOR2_X1   g784(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n986_));
  AND2_X1   g785(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n987_));
  NOR4_X1   g786(.A1(new_n979_), .A2(new_n342_), .A3(new_n986_), .A4(new_n987_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n986_), .B1(new_n979_), .B2(new_n342_), .ZN(new_n989_));
  OR2_X1    g788(.A1(new_n989_), .A2(KEYINPUT127), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n989_), .A2(KEYINPUT127), .ZN(new_n991_));
  AOI21_X1  g790(.A(new_n988_), .B1(new_n990_), .B2(new_n991_), .ZN(G1354gat));
  INV_X1    g791(.A(G218gat), .ZN(new_n993_));
  NOR3_X1   g792(.A1(new_n979_), .A2(new_n993_), .A3(new_n288_), .ZN(new_n994_));
  NAND3_X1  g793(.A1(new_n978_), .A2(new_n687_), .A3(new_n952_), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n994_), .B1(new_n993_), .B2(new_n995_), .ZN(G1355gat));
endmodule


