//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(G120gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT85), .B(G113gat), .Z(new_n206_));
  OR3_X1    g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G227gat), .A2(G233gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n209_), .B(new_n210_), .Z(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT30), .B(G15gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT31), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n211_), .B(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT26), .B1(new_n219_), .B2(KEYINPUT82), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT82), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(G190gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n220_), .B(new_n223_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  AND3_X1   g028(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n218_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n233_));
  INV_X1    g032(.A(new_n217_), .ZN(new_n234_));
  INV_X1    g033(.A(G183gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n219_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G176gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n229_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n238_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n232_), .A2(new_n233_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n233_), .B1(new_n232_), .B2(new_n246_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G71gat), .B(G99gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G43gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n249_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n214_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n214_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G233gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT86), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(KEYINPUT86), .ZN(new_n260_));
  OAI21_X1  g059(.A(G228gat), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT3), .Z(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT2), .Z(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n263_), .B1(new_n262_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n270_), .B2(new_n262_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n265_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n267_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(G211gat), .A2(G218gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G211gat), .A2(G218gat), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G197gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G204gat), .ZN(new_n283_));
  INV_X1    g082(.A(G204gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G197gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT21), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT87), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(G197gat), .B2(new_n284_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n284_), .A2(G197gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n288_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n281_), .B(new_n287_), .C1(new_n292_), .C2(KEYINPUT21), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n278_), .A2(KEYINPUT21), .A3(new_n279_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n292_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n293_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n261_), .B1(new_n277_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n261_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n275_), .B2(KEYINPUT29), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G78gat), .B(G106gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n275_), .A2(KEYINPUT29), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT28), .ZN(new_n307_));
  XOR2_X1   g106(.A(G22gat), .B(G50gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n275_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n209_), .A2(new_n275_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT4), .A3(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(KEYINPUT4), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n311_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n313_), .A2(new_n314_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n311_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G1gat), .B(G29gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT93), .B(G85gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT0), .B(G57gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n317_), .A2(new_n320_), .A3(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n282_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT87), .B1(new_n282_), .B2(G204gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n283_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT88), .B1(new_n335_), .B2(new_n294_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n292_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n280_), .B1(KEYINPUT21), .B2(new_n286_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n336_), .A2(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n225_), .A2(new_n224_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G190gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n245_), .A2(new_n242_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n345_), .A2(new_n218_), .B1(new_n346_), .B2(new_n238_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n232_), .A2(new_n246_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT84), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n232_), .A2(new_n233_), .A3(new_n246_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n341_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT20), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n348_), .B1(new_n353_), .B2(KEYINPUT90), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT90), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n355_), .A3(KEYINPUT20), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n332_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  AOI211_X1 g157(.A(new_n358_), .B(new_n331_), .C1(new_n341_), .C2(new_n347_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n299_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n357_), .A2(KEYINPUT94), .A3(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(KEYINPUT97), .ZN(new_n369_));
  XOR2_X1   g168(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n360_), .B1(new_n372_), .B2(KEYINPUT96), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n345_), .A2(new_n218_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n246_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n370_), .B1(new_n299_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT96), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n369_), .B(new_n331_), .C1(new_n373_), .C2(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n299_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT90), .B1(new_n380_), .B2(new_n358_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n348_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n381_), .A2(new_n332_), .A3(new_n356_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n377_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n372_), .A2(KEYINPUT96), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n360_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n369_), .B1(new_n387_), .B2(new_n331_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n363_), .A2(KEYINPUT32), .A3(new_n368_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n357_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(KEYINPUT94), .A3(new_n361_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n393_));
  INV_X1    g192(.A(new_n368_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n329_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n328_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT33), .B(new_n326_), .C1(new_n317_), .C2(new_n320_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n315_), .A2(new_n316_), .A3(new_n311_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n318_), .A2(new_n319_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n325_), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n391_), .A2(new_n404_), .A3(new_n368_), .A4(new_n361_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n394_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n352_), .A2(new_n355_), .A3(KEYINPUT20), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n355_), .B1(new_n352_), .B2(KEYINPUT20), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n348_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n368_), .B(new_n361_), .C1(new_n409_), .C2(new_n332_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n410_), .A3(KEYINPUT92), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n403_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n310_), .B1(new_n396_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n394_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT98), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n410_), .B2(KEYINPUT99), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT99), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n391_), .A2(new_n418_), .A3(new_n368_), .A4(new_n361_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT98), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n394_), .C1(new_n384_), .C2(new_n388_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n415_), .A2(new_n417_), .A3(new_n419_), .A4(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n310_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n411_), .A2(new_n416_), .A3(new_n405_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n329_), .A4(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n257_), .B1(new_n413_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n310_), .A3(new_n424_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT100), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT100), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n422_), .A2(new_n429_), .A3(new_n310_), .A4(new_n424_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n256_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n426_), .B1(new_n431_), .B2(new_n329_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G229gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT77), .B(G15gat), .ZN(new_n434_));
  INV_X1    g233(.A(G22gat), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n435_), .ZN(new_n437_));
  INV_X1    g236(.A(G1gat), .ZN(new_n438_));
  INV_X1    g237(.A(G8gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT14), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G1gat), .B(G8gat), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n442_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G43gat), .B(G50gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT71), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n446_), .A2(new_n447_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G29gat), .B(G36gat), .Z(new_n450_));
  OR3_X1    g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n445_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n453_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n433_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n453_), .B(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n454_), .B1(new_n459_), .B2(new_n445_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n457_), .B1(new_n460_), .B2(new_n433_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G169gat), .B(G197gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT81), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n461_), .B(new_n465_), .Z(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT69), .B(G71gat), .ZN(new_n467_));
  INV_X1    g266(.A(G78gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G64gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(KEYINPUT11), .A3(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(KEYINPUT11), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n469_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT67), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT7), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n478_));
  OAI22_X1  g277(.A1(new_n477_), .A2(new_n478_), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(KEYINPUT68), .A3(new_n481_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G85gat), .B(G92gat), .Z(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(KEYINPUT8), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT9), .ZN(new_n496_));
  INV_X1    g295(.A(G85gat), .ZN(new_n497_));
  INV_X1    g296(.A(G92gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT66), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n501_), .B(new_n502_), .C1(new_n491_), .C2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT10), .B(G99gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT65), .B(G106gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n488_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n494_), .A2(new_n495_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n492_), .A2(new_n493_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n493_), .B1(new_n492_), .B2(new_n508_), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT12), .B(new_n474_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT64), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n492_), .A2(new_n508_), .A3(new_n473_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT12), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n473_), .B1(new_n492_), .B2(new_n508_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n515_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n514_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G120gat), .B(G148gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(new_n284_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT5), .B(G176gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  NAND3_X1  g326(.A1(new_n520_), .A2(new_n523_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT13), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(KEYINPUT13), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n432_), .A2(new_n466_), .A3(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G190gat), .B(G218gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT36), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n492_), .A2(new_n508_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(new_n453_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(KEYINPUT70), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n509_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n544_), .B2(new_n459_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT75), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT75), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n544_), .A2(new_n459_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT73), .B(new_n549_), .C1(new_n557_), .C2(new_n542_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n540_), .B1(new_n562_), .B2(KEYINPUT76), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n553_), .A2(new_n555_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT76), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n538_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT74), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n563_), .A2(new_n566_), .B1(new_n564_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT78), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n445_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(new_n473_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577_));
  INV_X1    g376(.A(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT16), .B(G183gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n581_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n574_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n570_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n535_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n589_), .B2(new_n329_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT103), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n562_), .A2(new_n539_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n564_), .A2(new_n569_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(KEYINPUT37), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n570_), .B2(KEYINPUT37), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(new_n587_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n535_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n329_), .B(KEYINPUT101), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n597_), .A2(G1gat), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n591_), .A2(new_n602_), .ZN(G1324gat));
  INV_X1    g402(.A(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n422_), .A2(new_n424_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n439_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607_));
  INV_X1    g406(.A(new_n589_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n605_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n609_), .B2(G8gat), .ZN(new_n610_));
  AOI211_X1 g409(.A(KEYINPUT39), .B(new_n439_), .C1(new_n608_), .C2(new_n605_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT40), .B(new_n606_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1325gat));
  OAI21_X1  g415(.A(G15gat), .B1(new_n589_), .B2(new_n256_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n597_), .A2(G15gat), .A3(new_n256_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n589_), .B2(new_n310_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT42), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n604_), .A2(new_n435_), .A3(new_n423_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1327gat));
  NAND2_X1  g425(.A1(new_n428_), .A2(new_n430_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n329_), .A3(new_n257_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n426_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n534_), .A2(new_n466_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n539_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n562_), .A2(KEYINPUT76), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n593_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n586_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT106), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n630_), .A2(new_n638_), .A3(new_n631_), .A4(new_n635_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n329_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n534_), .A2(new_n466_), .A3(new_n586_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n630_), .A2(new_n644_), .A3(new_n645_), .A4(new_n595_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n592_), .A2(new_n593_), .A3(KEYINPUT37), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n634_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n432_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n644_), .B1(new_n652_), .B2(new_n645_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n643_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(G29gat), .A3(new_n598_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n641_), .B(new_n256_), .C1(new_n428_), .C2(new_n430_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n645_), .B(new_n595_), .C1(new_n658_), .C2(new_n426_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n650_), .A3(new_n646_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n643_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n642_), .B1(new_n657_), .B2(new_n662_), .ZN(G1328gat));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664_));
  INV_X1    g463(.A(G36gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n605_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n665_), .B1(new_n667_), .B2(new_n662_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n605_), .A2(KEYINPUT107), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n605_), .A2(KEYINPUT107), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n637_), .A2(new_n665_), .A3(new_n639_), .A4(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n664_), .B1(new_n668_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n672_), .B(KEYINPUT45), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n643_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT44), .B1(new_n661_), .B2(new_n643_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n666_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT46), .B(new_n676_), .C1(new_n679_), .C2(new_n665_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(new_n680_), .ZN(G1329gat));
  INV_X1    g480(.A(G43gat), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n256_), .A2(new_n682_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n656_), .A2(new_n662_), .A3(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n637_), .A2(new_n257_), .A3(new_n639_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n682_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(new_n682_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT47), .B1(new_n684_), .B2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n656_), .A2(new_n662_), .A3(new_n683_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n691_), .B(new_n692_), .C1(new_n688_), .C2(new_n687_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n640_), .B2(new_n423_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n656_), .A2(G50gat), .A3(new_n423_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g496(.A(new_n466_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n534_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n432_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n596_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n598_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n700_), .A2(G57gat), .A3(new_n641_), .A4(new_n588_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT109), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT109), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n703_), .A2(new_n705_), .A3(new_n706_), .ZN(G1332gat));
  NAND2_X1  g506(.A1(new_n700_), .A2(new_n588_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n671_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G64gat), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT48), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(G64gat), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT110), .Z(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n701_), .B2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n708_), .B2(new_n256_), .ZN(new_n715_));
  XOR2_X1   g514(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n256_), .A2(G71gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n701_), .B2(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n708_), .B2(new_n310_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n310_), .A2(G78gat), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT112), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n701_), .B2(new_n723_), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n700_), .A2(new_n635_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(KEYINPUT113), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n700_), .B2(new_n635_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n497_), .B1(new_n729_), .B2(new_n599_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n534_), .A2(new_n466_), .A3(new_n587_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT114), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n661_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n641_), .A2(G85gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT115), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n730_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(KEYINPUT116), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1336gat));
  NOR3_X1   g541(.A1(new_n733_), .A2(new_n498_), .A3(new_n709_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n725_), .B(KEYINPUT113), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n605_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n745_), .B2(new_n498_), .ZN(G1337gat));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n505_), .A3(new_n257_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G99gat), .B1(new_n733_), .B2(new_n256_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(new_n751_), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n661_), .A2(new_n423_), .A3(new_n732_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(G106gat), .A3(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n506_), .B(new_n423_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT53), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n759_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n757_), .A4(new_n756_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(G1339gat));
  NAND2_X1  g563(.A1(new_n461_), .A2(new_n465_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n455_), .A2(new_n456_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n465_), .B1(new_n766_), .B2(new_n433_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n460_), .A2(G229gat), .A3(G233gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(new_n528_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n512_), .A2(new_n519_), .A3(new_n771_), .A4(new_n514_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n527_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n474_), .A2(KEYINPUT12), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n543_), .B2(new_n509_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n517_), .B1(KEYINPUT12), .B2(new_n515_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n522_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n520_), .A2(new_n778_), .A3(KEYINPUT55), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n780_), .B2(KEYINPUT118), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n520_), .A2(new_n778_), .A3(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n772_), .A2(new_n773_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n779_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n781_), .A2(new_n788_), .A3(KEYINPUT119), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT119), .B1(new_n781_), .B2(new_n788_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(KEYINPUT58), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT120), .B1(new_n791_), .B2(new_n649_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n781_), .A2(new_n788_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n781_), .A2(new_n788_), .A3(KEYINPUT119), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n595_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n781_), .A2(new_n788_), .A3(KEYINPUT58), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n785_), .A2(new_n787_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n698_), .A3(new_n528_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n765_), .A2(new_n769_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n531_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n634_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(KEYINPUT57), .A3(new_n634_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n586_), .B1(new_n802_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n534_), .A2(new_n698_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n596_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n649_), .A2(new_n586_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n815_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n813_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n431_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n599_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826_), .B2(new_n698_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n822_), .A2(KEYINPUT59), .A3(new_n825_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  INV_X1    g628(.A(new_n801_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n595_), .A2(new_n798_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(KEYINPUT120), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n811_), .B1(new_n832_), .B2(new_n800_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n820_), .B1(new_n833_), .B2(new_n586_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n829_), .B1(new_n834_), .B2(new_n824_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n828_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n698_), .A2(G113gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT121), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n827_), .B1(new_n836_), .B2(new_n838_), .ZN(G1340gat));
  OAI21_X1  g638(.A(new_n203_), .B1(new_n699_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n826_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n203_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n828_), .A2(new_n835_), .A3(new_n699_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n203_), .ZN(G1341gat));
  AOI21_X1  g642(.A(G127gat), .B1(new_n826_), .B2(new_n586_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(G127gat), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n586_), .A2(KEYINPUT122), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(G127gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n844_), .B1(new_n836_), .B2(new_n848_), .ZN(G1342gat));
  NAND3_X1  g648(.A1(new_n834_), .A2(new_n570_), .A3(new_n824_), .ZN(new_n850_));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(KEYINPUT123), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n595_), .A2(G134gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT124), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n854_), .A2(new_n855_), .B1(new_n836_), .B2(new_n857_), .ZN(G1343gat));
  NOR3_X1   g657(.A1(new_n599_), .A2(new_n310_), .A3(new_n257_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n709_), .A2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT125), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n834_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n698_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n534_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n586_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n862_), .B2(new_n570_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n595_), .A2(G162gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT126), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n862_), .B2(new_n872_), .ZN(G1347gat));
  NOR3_X1   g672(.A1(new_n598_), .A2(new_n423_), .A3(new_n256_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n834_), .A2(new_n671_), .A3(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G169gat), .B1(new_n875_), .B2(new_n466_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n875_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n879_), .B(new_n698_), .C1(new_n241_), .C2(new_n240_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT62), .B(G169gat), .C1(new_n875_), .C2(new_n466_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  NOR2_X1   g681(.A1(new_n875_), .A2(new_n699_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n239_), .ZN(G1349gat));
  NAND3_X1  g683(.A1(new_n879_), .A2(new_n343_), .A3(new_n586_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G183gat), .B1(new_n875_), .B2(new_n587_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n875_), .B2(new_n649_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n570_), .A2(new_n344_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n875_), .B2(new_n889_), .ZN(G1351gat));
  NOR3_X1   g689(.A1(new_n257_), .A2(new_n641_), .A3(new_n310_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n671_), .B(new_n891_), .C1(new_n813_), .C2(new_n821_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n466_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n282_), .ZN(G1352gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n699_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n284_), .ZN(G1353gat));
  NOR2_X1   g695(.A1(new_n892_), .A2(new_n587_), .ZN(new_n897_));
  OR2_X1    g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT63), .B(G211gat), .Z(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n897_), .B2(new_n900_), .ZN(G1354gat));
  OAI21_X1  g700(.A(G218gat), .B1(new_n892_), .B2(new_n649_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n634_), .A2(G218gat), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n834_), .A2(new_n671_), .A3(new_n891_), .A4(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT127), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n902_), .A2(new_n907_), .A3(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1355gat));
endmodule


