//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_;
  XOR2_X1   g000(.A(G197gat), .B(G204gat), .Z(new_n202_));
  NAND3_X1  g001(.A1(new_n202_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT21), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n204_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n204_), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n209_), .A2(new_n202_), .A3(KEYINPUT89), .A4(KEYINPUT21), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT3), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n212_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n221_));
  OR2_X1    g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n222_), .B(new_n215_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n211_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G50gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n228_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G78gat), .B(G106gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G228gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(G22gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n231_), .A2(new_n234_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n235_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(G127gat), .A2(G134gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT87), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G127gat), .A2(G134gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n250_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n246_), .A2(new_n248_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT87), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n251_), .B1(new_n256_), .B2(new_n249_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(G227gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT81), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(KEYINPUT24), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267_));
  OR2_X1    g066(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(G190gat), .ZN(new_n271_));
  AND2_X1   g070(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT80), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n270_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277_));
  INV_X1    g076(.A(G183gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n279_), .A2(new_n280_), .B1(new_n267_), .B2(G190gat), .ZN(new_n281_));
  AND2_X1   g080(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT26), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT80), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n266_), .B1(new_n276_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT82), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT23), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(G183gat), .A3(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n290_), .A2(new_n292_), .B1(new_n293_), .B2(new_n264_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n266_), .B(KEYINPUT82), .C1(new_n276_), .C2(new_n285_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT22), .B(G169gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT83), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT84), .B(G176gat), .ZN(new_n299_));
  INV_X1    g098(.A(G169gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT83), .B1(new_n300_), .B2(KEYINPUT22), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n263_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT85), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n278_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n290_), .A2(new_n292_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(KEYINPUT85), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n296_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G71gat), .B(G99gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n310_), .B(KEYINPUT30), .ZN(new_n315_));
  INV_X1    g114(.A(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n261_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G15gat), .B(G43gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n314_), .A2(new_n317_), .A3(new_n261_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n323_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(new_n318_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n221_), .A2(new_n225_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n222_), .A2(KEYINPUT3), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n213_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n331_), .A2(new_n333_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n224_), .A3(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n336_), .C1(new_n254_), .C2(new_n257_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n252_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n256_), .A2(new_n251_), .A3(new_n249_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n338_), .B(new_n339_), .C1(new_n220_), .C2(new_n226_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n329_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n340_), .A3(KEYINPUT4), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n258_), .B(new_n344_), .C1(new_n226_), .C2(new_n220_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n342_), .B1(new_n346_), .B2(new_n328_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n347_), .B(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n324_), .A2(new_n327_), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT18), .B(G64gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G92gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n306_), .B1(G183gat), .B2(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n297_), .A2(new_n299_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n263_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT90), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT90), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n262_), .A2(new_n369_), .A3(KEYINPUT24), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n265_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n279_), .A2(new_n280_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n267_), .A2(G190gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n271_), .A3(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n294_), .A3(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n366_), .A2(new_n375_), .A3(KEYINPUT97), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT97), .B1(new_n366_), .B2(new_n375_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n211_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n310_), .B2(new_n211_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n363_), .B1(new_n379_), .B2(KEYINPUT20), .ZN(new_n380_));
  INV_X1    g179(.A(new_n211_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n296_), .A2(new_n309_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n366_), .A2(new_n375_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n211_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT91), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n211_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(KEYINPUT20), .A3(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(new_n362_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n360_), .B1(new_n380_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n362_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n310_), .A2(new_n211_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n211_), .A2(new_n383_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(KEYINPUT20), .A3(new_n363_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(KEYINPUT92), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n381_), .B1(new_n296_), .B2(new_n309_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n395_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n392_), .A2(new_n397_), .A3(new_n400_), .A4(new_n359_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n391_), .A2(KEYINPUT27), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n400_), .A3(new_n397_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n360_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT27), .B1(new_n404_), .B2(new_n401_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT100), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(KEYINPUT100), .ZN(new_n408_));
  AOI211_X1 g207(.A(new_n245_), .B(new_n355_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT99), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n380_), .B2(new_n390_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n347_), .B(new_n352_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n392_), .A2(new_n397_), .A3(new_n400_), .A4(new_n411_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n404_), .A2(new_n401_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT94), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n347_), .A2(new_n418_), .A3(KEYINPUT33), .A4(new_n352_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n328_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n420_));
  OAI211_X1 g219(.A(KEYINPUT33), .B(new_n352_), .C1(new_n420_), .C2(new_n341_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT94), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n352_), .B1(new_n420_), .B2(new_n341_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT95), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT95), .B(new_n352_), .C1(new_n420_), .C2(new_n341_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n343_), .A2(new_n345_), .A3(new_n328_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n337_), .A2(new_n340_), .A3(new_n329_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n353_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT96), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n423_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n416_), .B1(new_n417_), .B2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n435_), .A2(KEYINPUT98), .A3(new_n244_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT98), .B1(new_n435_), .B2(new_n244_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n354_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n402_), .A2(new_n405_), .A3(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n324_), .A2(new_n327_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n410_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n435_), .A2(new_n244_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n435_), .A2(KEYINPUT98), .A3(new_n244_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n439_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n441_), .A3(KEYINPUT99), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n409_), .B1(new_n443_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G57gat), .B(G64gat), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n452_), .A2(KEYINPUT11), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(KEYINPUT11), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G71gat), .B(G78gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G231gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G8gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G15gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n237_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G15gat), .A2(G22gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G1gat), .A2(G8gat), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n465_), .A2(new_n466_), .B1(KEYINPUT14), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n463_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n460_), .B(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G127gat), .B(G155gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G183gat), .B(G211gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  AND2_X1   g274(.A1(new_n475_), .A2(KEYINPUT17), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(KEYINPUT73), .Z(new_n478_));
  NOR2_X1   g277(.A1(new_n470_), .A2(new_n476_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(KEYINPUT17), .B2(new_n475_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G230gat), .ZN(new_n482_));
  INV_X1    g281(.A(G233gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT6), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  OR3_X1    g286(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G85gat), .B(G92gat), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(KEYINPUT65), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n491_), .B(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT10), .B(G99gat), .Z(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT64), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(KEYINPUT9), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT9), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(G85gat), .A3(G92gat), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n500_), .A2(new_n486_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n495_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(new_n458_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT12), .ZN(new_n507_));
  INV_X1    g306(.A(new_n505_), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n508_), .A2(KEYINPUT12), .A3(new_n458_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n484_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n506_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G120gat), .B(G148gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G204gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT5), .ZN(new_n515_));
  INV_X1    g314(.A(G176gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(KEYINPUT66), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT13), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT75), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G29gat), .B(G36gat), .ZN(new_n525_));
  INV_X1    g324(.A(G43gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(G50gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT68), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(G50gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n524_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n527_), .B(G50gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT68), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(KEYINPUT15), .A3(new_n531_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n469_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT76), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT76), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n535_), .B(KEYINPUT74), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n469_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n539_), .B(new_n540_), .C1(new_n538_), .C2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n542_), .B(new_n469_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n523_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT75), .B1(new_n545_), .B2(new_n546_), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT78), .B(G141gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G169gat), .B(G197gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT77), .B(G113gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n548_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n522_), .A2(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n451_), .A2(new_n481_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT34), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT35), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n508_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n505_), .A2(new_n535_), .B1(KEYINPUT35), .B2(new_n561_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n566_), .A2(KEYINPUT67), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT67), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n532_), .A2(new_n524_), .A3(new_n533_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT15), .B1(new_n536_), .B2(new_n531_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n505_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n567_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n565_), .B1(new_n568_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT67), .B1(new_n566_), .B2(new_n567_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n564_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(G134gat), .ZN(new_n580_));
  INV_X1    g379(.A(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n575_), .A2(KEYINPUT36), .A3(new_n578_), .A4(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n575_), .A2(new_n578_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT69), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n585_), .ZN(new_n589_));
  AOI211_X1 g388(.A(KEYINPUT69), .B(new_n589_), .C1(new_n575_), .C2(new_n578_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n584_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT37), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n584_), .B(new_n593_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n559_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT101), .ZN(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n414_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n591_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n559_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n354_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n601_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  NAND2_X1  g406(.A1(new_n407_), .A2(new_n408_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G8gat), .B1(new_n604_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT39), .ZN(new_n610_));
  INV_X1    g409(.A(G8gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n608_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n598_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g414(.A(G15gat), .B1(new_n604_), .B2(new_n441_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT41), .Z(new_n617_));
  NAND3_X1  g416(.A1(new_n598_), .A2(new_n464_), .A3(new_n442_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n604_), .B2(new_n244_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n598_), .A2(new_n237_), .A3(new_n245_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n409_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n449_), .A2(KEYINPUT99), .A3(new_n441_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT99), .B1(new_n449_), .B2(new_n441_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n481_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n558_), .A2(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n627_), .A2(new_n591_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n414_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n592_), .A2(KEYINPUT103), .A3(new_n594_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT103), .B1(new_n592_), .B2(new_n594_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT43), .B1(new_n451_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n595_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n451_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n627_), .A2(new_n640_), .A3(KEYINPUT104), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n635_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n629_), .B(KEYINPUT102), .Z(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n354_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n631_), .B1(new_n647_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g447(.A(G36gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n630_), .A2(new_n649_), .A3(new_n612_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n654_));
  AND3_X1   g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n646_), .A2(new_n608_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(new_n649_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n657_), .B(KEYINPUT46), .C1(new_n658_), .C2(new_n649_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1329gat));
  NAND2_X1  g462(.A1(new_n442_), .A2(G43gat), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n630_), .A2(new_n442_), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n646_), .A2(new_n664_), .B1(G43gat), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g466(.A1(new_n646_), .A2(KEYINPUT107), .A3(new_n244_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT107), .B1(new_n646_), .B2(new_n244_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(G50gat), .A3(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n630_), .A2(new_n230_), .A3(new_n245_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1331gat));
  INV_X1    g471(.A(new_n557_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n628_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n451_), .A2(new_n522_), .A3(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(new_n596_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G57gat), .B1(new_n676_), .B2(new_n414_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT108), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n603_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT109), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n414_), .A2(G57gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1332gat));
  INV_X1    g481(.A(G64gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n680_), .B2(new_n612_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT48), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n676_), .A2(new_n683_), .A3(new_n612_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1333gat));
  INV_X1    g486(.A(G71gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n680_), .B2(new_n442_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT49), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n676_), .A2(new_n688_), .A3(new_n442_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1334gat));
  INV_X1    g491(.A(G78gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n680_), .B2(new_n245_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT50), .Z(new_n695_));
  NAND3_X1  g494(.A1(new_n676_), .A2(new_n693_), .A3(new_n245_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1335gat));
  NOR3_X1   g496(.A1(new_n522_), .A2(new_n628_), .A3(new_n557_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n627_), .A2(new_n591_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G85gat), .B1(new_n699_), .B2(new_n414_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n642_), .A2(new_n698_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n414_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(new_n702_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g502(.A(G92gat), .B1(new_n699_), .B2(new_n612_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n701_), .A2(G92gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n612_), .ZN(G1337gat));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT51), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n701_), .A2(new_n442_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G99gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n699_), .A2(new_n496_), .A3(new_n442_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT110), .Z(new_n712_));
  AOI21_X1  g511(.A(new_n708_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n707_), .A2(KEYINPUT51), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n713_), .B(new_n714_), .Z(G1338gat));
  NAND3_X1  g514(.A1(new_n642_), .A2(new_n245_), .A3(new_n698_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n642_), .A2(KEYINPUT112), .A3(new_n245_), .A4(new_n698_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(G106gat), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT52), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n718_), .A2(new_n722_), .A3(G106gat), .A4(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n699_), .A2(new_n497_), .A3(new_n245_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n727_), .A3(new_n725_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1339gat));
  INV_X1    g530(.A(new_n522_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(new_n674_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n596_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT54), .Z(new_n735_));
  INV_X1    g534(.A(KEYINPUT118), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT55), .B1(new_n510_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n737_), .B1(new_n510_), .B2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n507_), .A2(new_n509_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n738_), .A2(new_n740_), .B1(new_n484_), .B2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n737_), .B(KEYINPUT55), .C1(new_n510_), .C2(new_n739_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n520_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n518_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT56), .B(new_n520_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n746_), .A2(new_n673_), .A3(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n539_), .B(new_n546_), .C1(new_n538_), .C2(new_n543_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n545_), .A2(new_n540_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n554_), .A3(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT116), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n555_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(KEYINPUT117), .A3(new_n521_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n555_), .A3(new_n521_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n603_), .B1(new_n748_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n736_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n760_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n744_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n744_), .A2(new_n745_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n764_), .A2(new_n557_), .A3(new_n518_), .A4(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n757_), .A3(new_n754_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n603_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n746_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n765_), .A3(new_n753_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n769_), .A2(KEYINPUT58), .A3(new_n765_), .A4(new_n753_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n595_), .A3(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n761_), .A2(new_n762_), .A3(new_n768_), .A4(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n735_), .B1(new_n775_), .B2(new_n481_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n612_), .A2(new_n354_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n442_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n776_), .A2(new_n245_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G113gat), .B1(new_n779_), .B2(new_n557_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n779_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NOR4_X1   g585(.A1(new_n776_), .A2(new_n245_), .A3(new_n778_), .A4(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n673_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n780_), .B1(new_n789_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g589(.A(G120gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n522_), .B2(KEYINPUT60), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n779_), .B(new_n792_), .C1(KEYINPUT60), .C2(new_n791_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n522_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n791_), .ZN(G1341gat));
  NOR2_X1   g594(.A1(new_n779_), .A2(new_n783_), .ZN(new_n796_));
  OAI211_X1 g595(.A(G127gat), .B(new_n628_), .C1(new_n796_), .C2(new_n787_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n776_), .A2(new_n481_), .A3(new_n245_), .A4(new_n778_), .ZN(new_n798_));
  OR3_X1    g597(.A1(new_n798_), .A2(KEYINPUT120), .A3(G127gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT120), .B1(new_n798_), .B2(G127gat), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n797_), .A2(new_n799_), .A3(new_n800_), .ZN(G1342gat));
  AOI21_X1  g600(.A(G134gat), .B1(new_n779_), .B2(new_n591_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n596_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g603(.A1(new_n775_), .A2(new_n481_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n735_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n442_), .A2(new_n244_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n777_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT121), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n673_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n522_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT122), .B(G148gat), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1345gat));
  NOR2_X1   g615(.A1(new_n811_), .A2(new_n481_), .ZN(new_n817_));
  XOR2_X1   g616(.A(KEYINPUT61), .B(G155gat), .Z(new_n818_));
  XNOR2_X1  g617(.A(new_n817_), .B(new_n818_), .ZN(G1346gat));
  NOR3_X1   g618(.A1(new_n811_), .A2(new_n581_), .A3(new_n634_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n581_), .B1(new_n811_), .B2(new_n603_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n821_), .A2(KEYINPUT123), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(KEYINPUT123), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n820_), .B1(new_n822_), .B2(new_n823_), .ZN(G1347gat));
  NOR2_X1   g623(.A1(new_n776_), .A2(new_n245_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n355_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n612_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G169gat), .B1(new_n827_), .B2(new_n673_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n557_), .A3(new_n297_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT62), .B(G169gat), .C1(new_n827_), .C2(new_n673_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n832_), .A3(new_n833_), .ZN(G1348gat));
  NOR3_X1   g633(.A1(new_n827_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n732_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n299_), .B2(new_n836_), .ZN(G1349gat));
  NAND4_X1  g636(.A1(new_n825_), .A2(new_n628_), .A3(new_n826_), .A4(new_n612_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n372_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n278_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT124), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n838_), .A2(new_n372_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n840_), .B1(new_n842_), .B2(new_n843_), .ZN(G1350gat));
  NAND4_X1  g643(.A1(new_n831_), .A2(new_n591_), .A3(new_n271_), .A4(new_n373_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n825_), .A2(new_n826_), .A3(new_n612_), .A4(new_n595_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n846_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT125), .B1(new_n846_), .B2(G190gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n847_), .B2(new_n848_), .ZN(G1351gat));
  NAND2_X1  g648(.A1(new_n612_), .A2(new_n808_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n776_), .A2(new_n414_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n557_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n732_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g654(.A(new_n850_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n807_), .A2(new_n354_), .A3(new_n628_), .A4(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT126), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n851_), .A2(new_n861_), .A3(new_n628_), .A4(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n860_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1354gat));
  NAND2_X1  g667(.A1(new_n851_), .A2(new_n591_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT127), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G218gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n851_), .A2(KEYINPUT127), .A3(new_n591_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n851_), .A2(G218gat), .A3(new_n595_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1355gat));
endmodule


