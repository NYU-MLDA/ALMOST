//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n968_, new_n969_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n977_, new_n978_, new_n979_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G120gat), .B(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT5), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G176gat), .B(G204gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT11), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G71gat), .B(G78gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n209_), .A2(KEYINPUT11), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n211_), .B1(KEYINPUT11), .B2(new_n209_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NOR3_X1   g021(.A1(KEYINPUT64), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n221_), .B(new_n222_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n226_), .A2(new_n224_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n218_), .B1(new_n225_), .B2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n217_), .B1(new_n231_), .B2(KEYINPUT67), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n233_), .B(new_n218_), .C1(new_n225_), .C2(new_n230_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n225_), .B2(new_n230_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT7), .ZN(new_n238_));
  AND3_X1   g037(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n238_), .A2(new_n241_), .A3(KEYINPUT65), .A4(new_n229_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n218_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n232_), .A2(new_n234_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT10), .B(G99gat), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n228_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n251_));
  INV_X1    g050(.A(G85gat), .ZN(new_n252_));
  INV_X1    g051(.A(G92gat), .ZN(new_n253_));
  OR3_X1    g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT9), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n250_), .A2(new_n251_), .A3(new_n254_), .A4(new_n241_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n216_), .B1(new_n248_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n216_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n234_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n238_), .A2(new_n241_), .A3(new_n229_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n233_), .B1(new_n260_), .B2(new_n218_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n259_), .A2(new_n261_), .A3(new_n217_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n246_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n258_), .B(new_n255_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n208_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  AOI211_X1 g067(.A(KEYINPUT68), .B(new_n266_), .C1(new_n257_), .C2(new_n264_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n257_), .A2(new_n264_), .A3(KEYINPUT12), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n231_), .A2(KEYINPUT67), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT8), .A3(new_n234_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n243_), .A2(new_n247_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n255_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n216_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n266_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n207_), .B1(new_n270_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n267_), .B1(new_n271_), .B2(new_n278_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n283_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT69), .B1(new_n284_), .B2(new_n207_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n258_), .B1(new_n275_), .B2(new_n255_), .ZN(new_n286_));
  AOI211_X1 g085(.A(new_n216_), .B(new_n256_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n267_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT68), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n265_), .A2(new_n208_), .A3(new_n267_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n292_));
  NOR4_X1   g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n283_), .A4(new_n206_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n282_), .B1(new_n285_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT13), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n280_), .A2(new_n290_), .A3(new_n289_), .A4(new_n207_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n292_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n270_), .A2(KEYINPUT69), .A3(new_n280_), .A4(new_n207_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n281_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT13), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G29gat), .B(G36gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G43gat), .B(G50gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n309_), .B(new_n312_), .Z(new_n313_));
  NAND2_X1  g112(.A1(G229gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n312_), .B(KEYINPUT15), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n309_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n309_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n312_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n318_), .A2(new_n320_), .A3(new_n314_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G113gat), .B(G141gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G169gat), .B(G197gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(KEYINPUT74), .A3(new_n328_), .ZN(new_n329_));
  OR3_X1    g128(.A1(new_n322_), .A2(KEYINPUT74), .A3(new_n325_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n303_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G231gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n309_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(new_n216_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT17), .ZN(new_n338_));
  XOR2_X1   g137(.A(G127gat), .B(G155gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT16), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G183gat), .B(G211gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  OR3_X1    g141(.A1(new_n337_), .A2(new_n338_), .A3(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(KEYINPUT17), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n333_), .A2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n349_));
  OAI21_X1  g148(.A(G169gat), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT79), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(G169gat), .C1(new_n348_), .C2(new_n349_), .ZN(new_n353_));
  INV_X1    g152(.A(G169gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(G176gat), .B1(new_n354_), .B2(KEYINPUT22), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G183gat), .ZN(new_n357_));
  INV_X1    g156(.A(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(KEYINPUT77), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT77), .B1(G183gat), .B2(G190gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n359_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n356_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n366_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n364_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n367_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n362_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n370_), .A2(KEYINPUT24), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n377_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n383_));
  OR3_X1    g182(.A1(new_n383_), .A2(new_n357_), .A3(KEYINPUT25), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT25), .B1(new_n383_), .B2(new_n357_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n376_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n371_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G15gat), .B(G43gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT31), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT81), .B(KEYINPUT82), .Z(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  XNOR2_X1  g198(.A(G113gat), .B(G120gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G127gat), .B(G134gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G134gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G127gat), .ZN(new_n406_));
  INV_X1    g205(.A(G127gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G134gat), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n406_), .A2(new_n408_), .A3(new_n403_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n401_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n408_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT83), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(new_n403_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n400_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n399_), .B(new_n415_), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n394_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT31), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n393_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n416_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G141gat), .A2(G148gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT84), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G141gat), .A2(G148gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n429_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n425_), .A2(new_n428_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n423_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(new_n426_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(KEYINPUT1), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G155gat), .A3(G162gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n441_), .A3(new_n433_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n415_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n432_), .A2(new_n435_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(new_n410_), .A3(KEYINPUT97), .A4(new_n414_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(KEYINPUT4), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n415_), .A2(new_n452_), .A3(new_n444_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(G85gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT0), .B(G57gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  NAND3_X1  g257(.A1(new_n446_), .A2(new_n450_), .A3(new_n448_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n454_), .B2(new_n459_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n422_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT95), .ZN(new_n467_));
  INV_X1    g266(.A(new_n370_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT77), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n367_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(KEYINPUT77), .A2(G183gat), .A3(G190gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT23), .A3(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n373_), .B2(new_n367_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n468_), .B1(new_n473_), .B2(new_n359_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n385_), .A2(new_n386_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n381_), .B1(new_n475_), .B2(new_n384_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n474_), .A2(new_n356_), .B1(new_n476_), .B2(new_n376_), .ZN(new_n477_));
  INV_X1    g276(.A(G211gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(G218gat), .ZN(new_n479_));
  INV_X1    g278(.A(G218gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(G211gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT89), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(G211gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(G218gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(G197gat), .A2(G204gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G197gat), .A2(G204gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT21), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n482_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT90), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n482_), .A2(new_n490_), .A3(new_n493_), .A4(new_n486_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n487_), .A2(new_n488_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(KEYINPUT21), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n482_), .A2(new_n486_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n492_), .A2(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n467_), .B1(new_n477_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n494_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(KEYINPUT95), .A3(new_n389_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT25), .B(G183gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n381_), .B1(new_n385_), .B2(new_n506_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n372_), .A2(new_n364_), .B1(G183gat), .B2(G190gat), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT23), .B1(new_n470_), .B2(new_n471_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n359_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT22), .B(G169gat), .ZN(new_n511_));
  INV_X1    g310(.A(G176gat), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n468_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n507_), .A2(new_n473_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT20), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G226gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT19), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n505_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n501_), .A2(new_n371_), .A3(new_n502_), .A4(new_n388_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(KEYINPUT20), .C1(new_n499_), .C2(new_n514_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n523_), .A2(KEYINPUT94), .A3(new_n519_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT94), .B1(new_n523_), .B2(new_n519_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G8gat), .B(G36gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT18), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G64gat), .B(G92gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT20), .B1(new_n499_), .B2(new_n514_), .ZN(new_n533_));
  AND4_X1   g332(.A1(new_n501_), .A2(new_n502_), .A3(new_n371_), .A4(new_n388_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n519_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT94), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n523_), .A2(KEYINPUT94), .A3(new_n519_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n539_), .A2(KEYINPUT96), .A3(new_n530_), .A4(new_n521_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n532_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n516_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n537_), .A2(new_n538_), .B1(new_n542_), .B2(new_n520_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT96), .B1(new_n543_), .B2(new_n530_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n466_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n530_), .B(new_n521_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n520_), .B1(new_n505_), .B2(new_n517_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n523_), .A2(new_n519_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n531_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n546_), .A2(KEYINPUT27), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G22gat), .B(G50gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n447_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n554_), .B1(new_n447_), .B2(new_n555_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n553_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n556_), .A3(new_n552_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n444_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n447_), .B2(new_n555_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n503_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT86), .B(G228gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT87), .B(G233gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G78gat), .B(G106gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT92), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n571_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT88), .Z(new_n577_));
  AND3_X1   g376(.A1(new_n444_), .A2(KEYINPUT85), .A3(KEYINPUT29), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT85), .B1(new_n444_), .B2(KEYINPUT29), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n503_), .B(new_n577_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n572_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n575_), .B1(new_n572_), .B2(new_n580_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n565_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n572_), .A2(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n574_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n572_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n564_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  AND4_X1   g387(.A1(KEYINPUT99), .A2(new_n545_), .A3(new_n551_), .A4(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n546_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n532_), .A3(new_n540_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n550_), .B1(new_n592_), .B2(new_n466_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT99), .B1(new_n593_), .B2(new_n588_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n465_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n583_), .A2(new_n587_), .A3(new_n463_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n550_), .A2(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n545_), .A2(KEYINPUT98), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT98), .B1(new_n545_), .B2(new_n597_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n588_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n449_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n458_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n446_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n460_), .A2(KEYINPUT33), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n454_), .A2(new_n606_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n591_), .A2(new_n532_), .A3(new_n608_), .A4(new_n540_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n461_), .A2(new_n462_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n530_), .A2(KEYINPUT32), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n610_), .B(new_n612_), .C1(new_n526_), .C2(new_n611_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n600_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n598_), .A2(new_n599_), .A3(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n595_), .B1(new_n615_), .B2(new_n422_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT71), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT36), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT70), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n276_), .A2(new_n623_), .A3(new_n317_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n256_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n317_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT70), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT34), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n625_), .A2(new_n312_), .B1(new_n632_), .B2(new_n631_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n628_), .B2(new_n635_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n622_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n623_), .B1(new_n276_), .B2(new_n317_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n625_), .A2(new_n626_), .A3(KEYINPUT70), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n633_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n621_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n646_), .A3(new_n636_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n639_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n347_), .A2(new_n616_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n202_), .B1(new_n650_), .B2(new_n610_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n643_), .A2(new_n646_), .A3(new_n636_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n622_), .B(KEYINPUT72), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n643_), .B2(new_n636_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT37), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT37), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n639_), .A2(new_n647_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n346_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n303_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT73), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n545_), .A2(new_n597_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n614_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n545_), .A2(new_n597_), .A3(KEYINPUT98), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n422_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n545_), .A2(new_n551_), .A3(new_n588_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n593_), .A2(KEYINPUT99), .A3(new_n588_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n464_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n665_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n331_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n660_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n202_), .A3(new_n610_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n651_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n675_), .B2(new_n674_), .ZN(G1324gat));
  INV_X1    g476(.A(new_n593_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n673_), .A2(new_n305_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n649_), .B2(new_n593_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n682_), .A2(G8gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n650_), .A2(KEYINPUT100), .A3(new_n678_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n680_), .A2(new_n684_), .A3(G8gat), .A4(new_n682_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n679_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT40), .B(new_n679_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1325gat));
  INV_X1    g490(.A(G15gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n673_), .A2(new_n692_), .A3(new_n422_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT101), .Z(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n650_), .B2(new_n422_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(new_n697_), .A3(new_n698_), .ZN(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n649_), .B2(new_n588_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  INV_X1    g500(.A(G22gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n673_), .A2(new_n702_), .A3(new_n600_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n655_), .A2(new_n657_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT102), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n665_), .B2(new_n670_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(KEYINPUT43), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n708_), .A2(KEYINPUT43), .B1(new_n616_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n346_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n333_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n705_), .B1(new_n710_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n616_), .B2(new_n707_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n709_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n665_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n595_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n712_), .C1(new_n716_), .C2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n714_), .A2(new_n610_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G29gat), .ZN(new_n722_));
  INV_X1    g521(.A(new_n648_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n346_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n302_), .A2(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n671_), .A2(new_n331_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n463_), .A2(G29gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n722_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n714_), .A2(new_n678_), .A3(new_n720_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT103), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n714_), .A2(new_n732_), .A3(new_n720_), .A4(new_n678_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n731_), .A2(G36gat), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G36gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n735_), .A3(new_n678_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT45), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n734_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1329gat));
  AND2_X1   g542(.A1(new_n422_), .A2(G43gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n714_), .A2(new_n720_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n714_), .A2(KEYINPUT105), .A3(new_n720_), .A4(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G43gat), .B1(new_n726_), .B2(new_n422_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT106), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT47), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n749_), .A2(new_n751_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1330gat));
  OR3_X1    g555(.A1(new_n727_), .A2(G50gat), .A3(new_n588_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n714_), .A2(new_n600_), .A3(new_n720_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n758_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT107), .B1(new_n758_), .B2(G50gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G1331gat));
  NAND2_X1  g560(.A1(new_n302_), .A2(new_n658_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT108), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n616_), .A3(new_n331_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT109), .Z(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n610_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n303_), .A2(new_n332_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n616_), .A2(new_n711_), .A3(new_n648_), .A4(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT110), .Z(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n610_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n766_), .B2(new_n771_), .ZN(G1332gat));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n773_), .A3(new_n678_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n678_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G64gat), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT48), .B(new_n773_), .C1(new_n770_), .C2(new_n678_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n765_), .A2(new_n780_), .A3(new_n422_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n770_), .A2(new_n422_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G71gat), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT49), .B(new_n780_), .C1(new_n770_), .C2(new_n422_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1334gat));
  INV_X1    g585(.A(G78gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n765_), .A2(new_n787_), .A3(new_n600_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n770_), .A2(new_n600_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G78gat), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT50), .B(new_n787_), .C1(new_n770_), .C2(new_n600_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(G1335gat));
  NOR4_X1   g592(.A1(new_n671_), .A2(new_n332_), .A3(new_n303_), .A4(new_n724_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n252_), .A3(new_n610_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n768_), .A2(new_n346_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n710_), .A2(new_n463_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n252_), .ZN(G1336gat));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n253_), .A3(new_n678_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n710_), .A2(new_n593_), .A3(new_n796_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n253_), .ZN(G1337gat));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n422_), .A3(new_n249_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n710_), .A2(new_n796_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n422_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n804_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT111), .B1(new_n804_), .B2(G99gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT51), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n802_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1338gat));
  NAND3_X1  g610(.A1(new_n794_), .A2(new_n228_), .A3(new_n600_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n803_), .A2(new_n600_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n813_), .A2(G106gat), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n813_), .B2(G106gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n812_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT53), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n812_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1339gat));
  NAND4_X1  g620(.A1(new_n296_), .A2(new_n658_), .A3(new_n331_), .A4(new_n301_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT54), .B1(new_n822_), .B2(KEYINPUT113), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825_));
  INV_X1    g624(.A(new_n822_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n822_), .A2(KEYINPUT113), .A3(KEYINPUT114), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n826_), .A2(new_n827_), .A3(new_n825_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT114), .B1(new_n822_), .B2(KEYINPUT113), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n823_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n313_), .A2(new_n314_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n318_), .A2(new_n320_), .A3(new_n315_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n327_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n326_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n280_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT55), .B1(new_n283_), .B2(KEYINPUT115), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n279_), .B2(new_n266_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n271_), .A2(KEYINPUT116), .A3(new_n267_), .A4(new_n278_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n842_), .A2(new_n843_), .A3(new_n845_), .A4(new_n846_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n206_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n206_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n839_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n706_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT58), .B(new_n839_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n838_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n294_), .A2(KEYINPUT118), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n300_), .B2(new_n838_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n331_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT117), .B(new_n863_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n648_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(KEYINPUT57), .A3(new_n648_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n857_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n834_), .B1(new_n873_), .B2(new_n346_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n668_), .A2(new_n669_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n610_), .A3(new_n422_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n874_), .B2(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n830_), .A2(new_n833_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n868_), .A2(KEYINPUT57), .A3(new_n648_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n870_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n868_), .B2(new_n648_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n852_), .A2(new_n854_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n879_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n878_), .B1(new_n883_), .B2(new_n711_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n876_), .A2(KEYINPUT59), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n877_), .A2(new_n886_), .A3(new_n332_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G113gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n874_), .A2(new_n876_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n331_), .A2(G113gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n888_), .B1(new_n890_), .B2(new_n891_), .ZN(G1340gat));
  NAND3_X1  g691(.A1(new_n877_), .A2(new_n886_), .A3(new_n302_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G120gat), .ZN(new_n894_));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n303_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(KEYINPUT60), .B2(new_n895_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n894_), .B1(new_n890_), .B2(new_n897_), .ZN(G1341gat));
  AOI21_X1  g697(.A(G127gat), .B1(new_n889_), .B2(new_n711_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n877_), .A2(new_n886_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n346_), .A2(new_n407_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT121), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n900_), .B2(new_n902_), .ZN(G1342gat));
  INV_X1    g702(.A(new_n706_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n877_), .A2(new_n886_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G134gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n889_), .A2(new_n405_), .A3(new_n723_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1343gat));
  NOR4_X1   g707(.A1(new_n678_), .A2(new_n422_), .A3(new_n588_), .A4(new_n463_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n859_), .A2(new_n861_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n865_), .B2(new_n864_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n723_), .B1(new_n912_), .B2(new_n867_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n872_), .B1(new_n913_), .B2(new_n880_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n855_), .A2(new_n856_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n346_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n910_), .B1(new_n916_), .B2(new_n878_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n332_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n917_), .B2(new_n302_), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n874_), .A2(KEYINPUT123), .A3(new_n303_), .A4(new_n910_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(G148gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n921_), .A2(new_n922_), .A3(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n879_), .A2(new_n881_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n711_), .B1(new_n926_), .B2(new_n857_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n302_), .B(new_n909_), .C1(new_n927_), .C2(new_n834_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT123), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n917_), .A2(new_n920_), .A3(new_n302_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n923_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n925_), .A2(new_n931_), .ZN(G1345gat));
  NAND2_X1  g731(.A1(new_n917_), .A2(new_n711_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT61), .B(G155gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1346gat));
  AND3_X1   g734(.A1(new_n917_), .A2(G162gat), .A3(new_n707_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n874_), .A2(new_n648_), .A3(new_n910_), .ZN(new_n937_));
  OR3_X1    g736(.A1(new_n937_), .A2(KEYINPUT124), .A3(G162gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT124), .B1(new_n937_), .B2(G162gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n936_), .B1(new_n938_), .B2(new_n939_), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n464_), .A2(new_n593_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n600_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n884_), .A2(new_n332_), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n945_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n511_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n948_), .B1(new_n944_), .B2(new_n354_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n946_), .A2(new_n947_), .A3(new_n949_), .ZN(G1348gat));
  AND2_X1   g749(.A1(new_n884_), .A2(new_n943_), .ZN(new_n951_));
  AOI21_X1  g750(.A(G176gat), .B1(new_n951_), .B2(new_n302_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n916_), .A2(new_n878_), .ZN(new_n953_));
  AOI21_X1  g752(.A(KEYINPUT125), .B1(new_n953_), .B2(new_n588_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n874_), .A2(new_n955_), .A3(new_n600_), .ZN(new_n956_));
  OR2_X1    g755(.A1(new_n954_), .A2(new_n956_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n942_), .A2(new_n303_), .A3(new_n512_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n952_), .B1(new_n957_), .B2(new_n958_), .ZN(G1349gat));
  NOR2_X1   g758(.A1(new_n346_), .A2(new_n506_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n884_), .A2(new_n943_), .A3(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(KEYINPUT126), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n884_), .A2(new_n963_), .A3(new_n943_), .A4(new_n960_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n711_), .B(new_n941_), .C1(new_n954_), .C2(new_n956_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n966_), .B2(new_n357_), .ZN(G1350gat));
  NAND3_X1  g766(.A1(new_n951_), .A2(new_n385_), .A3(new_n723_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n951_), .A2(new_n904_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n358_), .ZN(G1351gat));
  NOR4_X1   g769(.A1(new_n874_), .A2(new_n593_), .A3(new_n422_), .A4(new_n596_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(KEYINPUT127), .B(G197gat), .ZN(new_n972_));
  AND3_X1   g771(.A1(new_n971_), .A2(new_n332_), .A3(new_n972_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n972_), .B1(new_n971_), .B2(new_n332_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n973_), .A2(new_n974_), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n971_), .A2(new_n302_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(G204gat), .ZN(new_n977_));
  INV_X1    g776(.A(G204gat), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n971_), .A2(new_n978_), .A3(new_n302_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n977_), .A2(new_n979_), .ZN(G1353gat));
  OR2_X1    g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n971_), .B2(new_n711_), .ZN(new_n982_));
  AND2_X1   g781(.A1(new_n971_), .A2(new_n711_), .ZN(new_n983_));
  XOR2_X1   g782(.A(KEYINPUT63), .B(G211gat), .Z(new_n984_));
  AOI21_X1  g783(.A(new_n982_), .B1(new_n983_), .B2(new_n984_), .ZN(G1354gat));
  NAND3_X1  g784(.A1(new_n971_), .A2(new_n480_), .A3(new_n723_), .ZN(new_n986_));
  AND2_X1   g785(.A1(new_n971_), .A2(new_n904_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n986_), .B1(new_n987_), .B2(new_n480_), .ZN(G1355gat));
endmodule


