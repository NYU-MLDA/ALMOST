//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n207_), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT7), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT64), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n217_), .B1(new_n223_), .B2(new_n206_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n206_), .A2(new_n217_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(new_n212_), .B2(new_n221_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n230_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n227_), .B(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G230gat), .A3(G233gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT12), .B1(new_n227_), .B2(new_n234_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n227_), .A2(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n227_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT65), .B(new_n216_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(KEYINPUT12), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n240_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G120gat), .B(G148gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G176gat), .B(G204gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n236_), .A2(new_n247_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT13), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT13), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT69), .B(G15gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G22gat), .ZN(new_n265_));
  INV_X1    g064(.A(G8gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G1gat), .B(G8gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n265_), .A2(new_n271_), .A3(new_n267_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G29gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G43gat), .B(G50gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n273_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G229gat), .A2(G233gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT74), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n273_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n276_), .B(KEYINPUT15), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT75), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n270_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n273_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n283_), .A2(new_n278_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289_));
  INV_X1    g088(.A(new_n278_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n280_), .A2(new_n276_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n289_), .B(new_n290_), .C1(new_n291_), .C2(new_n284_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n279_), .A2(new_n288_), .A3(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G113gat), .B(G141gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(G169gat), .B(G197gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n279_), .A2(new_n288_), .A3(new_n292_), .A4(new_n296_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n263_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n234_), .ZN(new_n301_));
  INV_X1    g100(.A(G231gat), .ZN(new_n302_));
  INV_X1    g101(.A(G233gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n270_), .A2(new_n272_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n301_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n273_), .A2(new_n304_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n270_), .A2(new_n272_), .A3(new_n305_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n234_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G127gat), .B(G155gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT16), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G183gat), .B(G211gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT70), .B1(new_n312_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n321_));
  AOI211_X1 g120(.A(new_n321_), .B(new_n318_), .C1(new_n308_), .C2(new_n311_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n316_), .B(KEYINPUT17), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n308_), .A2(new_n311_), .A3(KEYINPUT71), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT71), .B1(new_n308_), .B2(new_n311_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n312_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n326_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT72), .B1(new_n334_), .B2(new_n325_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n324_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT73), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n329_), .A2(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(KEYINPUT72), .A3(new_n325_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n324_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n300_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n276_), .B(new_n216_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT35), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G232gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT34), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n346_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n242_), .A2(new_n281_), .A3(new_n243_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n350_), .A2(new_n347_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n351_), .B(new_n352_), .C1(new_n347_), .C2(new_n350_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G190gat), .B(G218gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G134gat), .B(G162gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT67), .B(KEYINPUT36), .Z(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n355_), .A2(new_n356_), .A3(new_n363_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT68), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n361_), .B(KEYINPUT36), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT31), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n380_), .B(new_n381_), .C1(G183gat), .C2(G190gat), .ZN(new_n382_));
  INV_X1    g181(.A(G176gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT79), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G176gat), .ZN(new_n386_));
  INV_X1    g185(.A(G169gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT22), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT22), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G169gat), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .A4(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n382_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT25), .B(G183gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398_));
  INV_X1    g197(.A(G190gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT26), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n399_), .A2(KEYINPUT26), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n397_), .B(new_n400_), .C1(new_n401_), .C2(new_n398_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n380_), .A2(new_n381_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT78), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n387_), .A3(new_n383_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n405_), .A2(KEYINPUT24), .A3(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n405_), .A2(new_n406_), .B1(KEYINPUT24), .B2(new_n393_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n402_), .B(new_n403_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n396_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT81), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n396_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G71gat), .B(G99gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT82), .B(G43gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n414_), .A2(new_n417_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G127gat), .B(G134gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n418_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n414_), .A2(new_n417_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n414_), .A2(new_n417_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n377_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n422_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n376_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G22gat), .B(G50gat), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G141gat), .A2(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n440_), .A2(KEYINPUT1), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(KEYINPUT1), .B2(new_n440_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n439_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(G155gat), .B(G162gat), .Z(new_n445_));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n436_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT2), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(G141gat), .B2(G148gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n438_), .A2(KEYINPUT2), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n453_));
  NOR3_X1   g252(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n446_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n445_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT84), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n458_), .B(new_n445_), .C1(new_n452_), .C2(new_n455_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n444_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT29), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n435_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n434_), .A3(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G211gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(G218gat), .ZN(new_n472_));
  INV_X1    g271(.A(G218gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(G211gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT88), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(G211gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(G218gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481_));
  INV_X1    g280(.A(G204gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(G197gat), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT21), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487_));
  INV_X1    g286(.A(G197gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(G204gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT87), .B1(new_n482_), .B2(G197gat), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n485_), .A2(new_n486_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n486_), .B1(G197gat), .B2(G204gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n483_), .A2(new_n484_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(G197gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n480_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n485_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n496_), .A2(KEYINPUT21), .A3(new_n479_), .A4(new_n475_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n499_));
  INV_X1    g298(.A(G228gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(new_n303_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  OAI221_X1 g301(.A(new_n498_), .B1(new_n500_), .B2(new_n303_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G78gat), .B(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n505_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n470_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n506_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n504_), .A2(new_n510_), .A3(new_n505_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n470_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT90), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n517_));
  AOI211_X1 g316(.A(new_n517_), .B(new_n470_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n509_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G8gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT18), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G64gat), .B(G92gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n413_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n412_), .B1(new_n396_), .B2(new_n409_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n498_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n382_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n407_), .A2(new_n408_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n397_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT26), .B(G190gat), .Z(new_n531_));
  OAI21_X1  g330(.A(new_n403_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n528_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n498_), .A2(KEYINPUT91), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT91), .B1(new_n498_), .B2(new_n533_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT20), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n527_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G226gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT19), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT20), .B1(new_n498_), .B2(new_n533_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT97), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n498_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT98), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n541_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n542_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n498_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n546_), .B(new_n539_), .C1(new_n549_), .C2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n524_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n539_), .B1(new_n527_), .B2(new_n536_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT20), .B(new_n540_), .C1(new_n498_), .C2(new_n533_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT92), .B1(new_n551_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n544_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n555_), .A2(new_n557_), .A3(new_n523_), .A4(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n561_), .A2(KEYINPUT27), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n524_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT27), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n554_), .A2(new_n562_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G1gat), .B(G29gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(G85gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT0), .B(G57gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n444_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n459_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n436_), .A2(new_n447_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT83), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n438_), .A2(KEYINPUT2), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n449_), .A2(G141gat), .A3(G148gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n575_), .A2(new_n578_), .A3(new_n453_), .A4(new_n448_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n458_), .B1(new_n579_), .B2(new_n445_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n572_), .B1(new_n573_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n422_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n457_), .A2(new_n459_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n572_), .A3(new_n424_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(KEYINPUT4), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G225gat), .A2(G233gat), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT4), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(new_n589_), .A3(new_n422_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT93), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n424_), .B1(new_n583_), .B2(new_n572_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT93), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n582_), .A2(new_n586_), .A3(new_n584_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n571_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n571_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n588_), .B2(new_n595_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n519_), .A2(new_n567_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n509_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n507_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n510_), .B2(new_n508_), .ZN(new_n605_));
  AOI211_X1 g404(.A(KEYINPUT89), .B(new_n507_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n515_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n517_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n514_), .A2(KEYINPUT90), .A3(new_n515_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n603_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n600_), .B2(KEYINPUT33), .ZN(new_n612_));
  INV_X1    g411(.A(new_n599_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n591_), .A2(new_n594_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n585_), .A2(new_n587_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(KEYINPUT94), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n613_), .B(KEYINPUT33), .C1(new_n614_), .C2(new_n615_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n564_), .A2(new_n561_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n444_), .B(new_n422_), .C1(new_n457_), .C2(new_n459_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n592_), .B2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n582_), .A2(KEYINPUT95), .A3(new_n584_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n587_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n571_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n626_), .A2(KEYINPUT96), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT96), .B1(new_n626_), .B2(new_n627_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n595_), .A2(new_n586_), .A3(new_n585_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n619_), .A2(new_n621_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n523_), .A2(KEYINPUT32), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI22_X1  g433(.A1(new_n598_), .A2(new_n600_), .B1(new_n563_), .B2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n539_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n636_), .A2(KEYINPUT98), .B1(new_n540_), .B2(new_n537_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n637_), .B2(new_n552_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n610_), .B1(new_n632_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n433_), .B1(new_n602_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n567_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n433_), .A2(new_n601_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n642_), .A2(new_n519_), .A3(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n344_), .B(new_n371_), .C1(new_n641_), .C2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT100), .Z(new_n646_));
  INV_X1    g445(.A(new_n601_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n202_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n341_), .B1(new_n340_), .B2(new_n324_), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT73), .B(new_n323_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n371_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n369_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT37), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n652_), .A2(new_n654_), .A3(new_n263_), .A4(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n602_), .A2(new_n640_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n644_), .B1(new_n658_), .B2(new_n432_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n299_), .B(KEYINPUT76), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT99), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n662_));
  INV_X1    g461(.A(new_n660_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n662_), .B(new_n663_), .C1(new_n641_), .C2(new_n644_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n657_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n202_), .A3(new_n647_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n648_), .B1(new_n649_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n649_), .B2(new_n666_), .ZN(G1324gat));
  OR3_X1    g467(.A1(new_n645_), .A2(KEYINPUT102), .A3(new_n567_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT102), .B1(new_n645_), .B2(new_n567_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(G8gat), .A3(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n567_), .A2(G8gat), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n665_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(KEYINPUT101), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n665_), .A2(KEYINPUT101), .A3(new_n675_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n673_), .B(new_n674_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n676_), .B(KEYINPUT101), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n683_), .A2(new_n673_), .A3(new_n674_), .A4(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1325gat));
  NAND2_X1  g484(.A1(new_n646_), .A2(new_n433_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G15gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n665_), .A2(new_n373_), .A3(new_n433_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n688_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n646_), .A2(new_n519_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G22gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n665_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n610_), .A2(G22gat), .ZN(new_n699_));
  OAI22_X1  g498(.A1(new_n696_), .A2(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n661_), .A2(new_n664_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n652_), .A2(new_n262_), .A3(new_n371_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G29gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n647_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n654_), .A2(new_n656_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n659_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n300_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT43), .B(new_n707_), .C1(new_n641_), .C2(new_n644_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n709_), .A2(new_n343_), .A3(new_n710_), .A4(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT107), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n712_), .A2(new_n713_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n601_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n705_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(G36gat), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n701_), .A2(new_n726_), .A3(new_n642_), .A4(new_n702_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT45), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n642_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n728_), .B1(new_n730_), .B2(new_n726_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n728_), .B(KEYINPUT46), .C1(new_n730_), .C2(new_n726_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1329gat));
  INV_X1    g534(.A(new_n720_), .ZN(new_n736_));
  INV_X1    g535(.A(G43gat), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n432_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n717_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n716_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n736_), .B(new_n738_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n703_), .A2(new_n433_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n737_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n741_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1330gat));
  AOI21_X1  g548(.A(G50gat), .B1(new_n703_), .B2(new_n519_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n720_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n519_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(G1331gat));
  INV_X1    g552(.A(G57gat), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n655_), .A2(KEYINPUT37), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n653_), .B(new_n369_), .C1(new_n364_), .C2(new_n366_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n343_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n262_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT110), .Z(new_n759_));
  NOR2_X1   g558(.A1(new_n659_), .A2(new_n299_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n754_), .B1(new_n761_), .B2(new_n601_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n659_), .A2(new_n655_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(new_n660_), .A3(new_n262_), .A4(new_n652_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n764_), .A2(new_n754_), .A3(new_n601_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(KEYINPUT111), .B2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(KEYINPUT111), .B2(new_n765_), .ZN(G1332gat));
  OAI21_X1  g566(.A(G64gat), .B1(new_n764_), .B2(new_n567_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT48), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n567_), .A2(G64gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n761_), .B2(new_n770_), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n764_), .B2(new_n432_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT49), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n432_), .A2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n761_), .B2(new_n774_), .ZN(G1334gat));
  OAI21_X1  g574(.A(G78gat), .B1(new_n764_), .B2(new_n610_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n610_), .A2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n761_), .B2(new_n779_), .ZN(G1335gat));
  OAI21_X1  g579(.A(new_n707_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n652_), .B1(new_n781_), .B2(new_n706_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n263_), .A2(new_n299_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n711_), .A3(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n601_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n760_), .A2(new_n262_), .A3(new_n343_), .A4(new_n655_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n213_), .A3(new_n647_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(G1336gat));
  OAI21_X1  g588(.A(G92gat), .B1(new_n784_), .B2(new_n567_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n214_), .A3(new_n642_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n784_), .B2(new_n432_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n433_), .A3(new_n203_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT113), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n795_), .B(new_n797_), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n787_), .A2(new_n204_), .A3(new_n519_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n782_), .A2(new_n519_), .A3(new_n711_), .A4(new_n783_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(G106gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(G106gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n757_), .A2(new_n806_), .A3(new_n660_), .A4(new_n263_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT54), .B1(new_n657_), .B2(new_n663_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n283_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT115), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n283_), .A2(new_n814_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n290_), .A3(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n277_), .A2(new_n290_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n296_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n298_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n811_), .B1(new_n820_), .B2(new_n258_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n257_), .A2(new_n819_), .A3(KEYINPUT116), .A4(new_n298_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n240_), .B1(new_n239_), .B2(new_n246_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n247_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n239_), .A2(new_n246_), .A3(KEYINPUT55), .A4(new_n240_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n255_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(new_n829_), .A3(KEYINPUT56), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n256_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n823_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n810_), .B1(new_n837_), .B2(new_n655_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n823_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n833_), .A2(new_n832_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n836_), .B1(new_n840_), .B2(new_n830_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n655_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT57), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n820_), .A2(new_n835_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n832_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n844_), .B(KEYINPUT58), .C1(new_n845_), .C2(new_n846_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n707_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n838_), .A2(new_n843_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n809_), .B1(new_n343_), .B2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n642_), .A2(new_n519_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n432_), .A2(new_n601_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n851_), .B1(new_n842_), .B2(KEYINPUT57), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n837_), .A2(new_n810_), .A3(new_n655_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n343_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT117), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n852_), .A2(new_n862_), .A3(new_n343_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n809_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n857_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866_), .B2(new_n660_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n809_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n860_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n856_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n299_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n872_), .A2(G113gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n867_), .B1(new_n871_), .B2(new_n873_), .ZN(G1340gat));
  OAI21_X1  g673(.A(G120gat), .B1(new_n866_), .B2(new_n263_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n876_));
  AOI21_X1  g675(.A(G120gat), .B1(new_n262_), .B2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT118), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n876_), .B2(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n877_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n875_), .B1(new_n871_), .B2(new_n881_), .ZN(G1341gat));
  INV_X1    g681(.A(G127gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n343_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n857_), .B(new_n884_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n871_), .B2(new_n343_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(KEYINPUT119), .A3(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n708_), .A2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n857_), .B(new_n893_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n871_), .B2(new_n371_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT120), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(new_n898_), .A3(new_n895_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n642_), .A2(new_n610_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n647_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n853_), .A2(new_n433_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n299_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n262_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g706(.A1(new_n869_), .A2(new_n647_), .A3(new_n432_), .A4(new_n901_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT121), .B1(new_n908_), .B2(new_n343_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n903_), .A2(new_n910_), .A3(new_n652_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT61), .B(G155gat), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n909_), .A2(new_n911_), .A3(new_n913_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1346gat));
  OR3_X1    g716(.A1(new_n908_), .A2(G162gat), .A3(new_n371_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G162gat), .B1(new_n908_), .B2(new_n708_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1347gat));
  INV_X1    g719(.A(new_n863_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n862_), .B1(new_n852_), .B2(new_n343_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n868_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n567_), .A2(new_n647_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n433_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n519_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927_), .B2(new_n872_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n926_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n861_), .A2(new_n863_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n868_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n933_), .A2(new_n388_), .A3(new_n390_), .A4(new_n299_), .ZN(new_n934_));
  OAI211_X1 g733(.A(KEYINPUT62), .B(G169gat), .C1(new_n927_), .C2(new_n872_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n930_), .A2(new_n934_), .A3(new_n935_), .ZN(G1348gat));
  NAND2_X1  g735(.A1(new_n869_), .A2(new_n610_), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n937_), .A2(new_n383_), .A3(new_n263_), .A4(new_n925_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n933_), .A2(new_n262_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT79), .B(G176gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(G1349gat));
  INV_X1    g740(.A(G183gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n652_), .A2(new_n433_), .A3(new_n924_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n937_), .B2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n652_), .A2(new_n530_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n927_), .B2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(KEYINPUT122), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n944_), .B(new_n948_), .C1(new_n927_), .C2(new_n945_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n927_), .B2(new_n708_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n371_), .A2(new_n531_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n933_), .A2(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n951_), .A2(KEYINPUT123), .A3(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n399_), .B1(new_n933_), .B2(new_n707_), .ZN(new_n956_));
  NOR4_X1   g755(.A1(new_n864_), .A2(new_n531_), .A3(new_n371_), .A4(new_n931_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n958_), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n853_), .A2(new_n433_), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n610_), .A2(new_n567_), .A3(new_n647_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n872_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(new_n488_), .ZN(G1352gat));
  NAND3_X1  g763(.A1(new_n960_), .A2(new_n262_), .A3(new_n961_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n966_), .B1(new_n482_), .B2(new_n965_), .ZN(G1353gat));
  NOR2_X1   g766(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(KEYINPUT125), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT126), .ZN(new_n970_));
  AND2_X1   g769(.A1(new_n960_), .A2(new_n961_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n343_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n972_));
  XOR2_X1   g771(.A(new_n972_), .B(KEYINPUT124), .Z(new_n973_));
  AOI21_X1  g772(.A(new_n970_), .B1(new_n971_), .B2(new_n973_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n971_), .A2(new_n973_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n969_), .A2(new_n976_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n974_), .B1(new_n975_), .B2(new_n977_), .ZN(G1354gat));
  NAND3_X1  g777(.A1(new_n971_), .A2(new_n473_), .A3(new_n655_), .ZN(new_n979_));
  OAI21_X1  g778(.A(G218gat), .B1(new_n962_), .B2(new_n708_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1355gat));
endmodule


