//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  OR2_X1    g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR3_X1   g007(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n206_), .B1(new_n210_), .B2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n203_), .B1(new_n216_), .B2(KEYINPUT67), .ZN(new_n217_));
  INV_X1    g016(.A(new_n206_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n212_), .A2(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n207_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n218_), .B1(new_n219_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n215_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT66), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n210_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n206_), .A2(KEYINPUT8), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n217_), .A2(new_n227_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n204_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n234_));
  OR2_X1    g033(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(G85gat), .A4(G92gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n204_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n205_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT10), .B(G99gat), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n222_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n229_), .A2(new_n230_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n202_), .B1(new_n233_), .B2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G29gat), .B(G36gat), .Z(new_n244_));
  XOR2_X1   g043(.A(G43gat), .B(G50gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT15), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n231_), .A2(new_n232_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT8), .B1(new_n225_), .B2(new_n226_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n216_), .A2(KEYINPUT67), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n242_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT68), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n243_), .A2(new_n247_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT73), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n217_), .A2(new_n227_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n242_), .B1(new_n260_), .B2(new_n248_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n261_), .B2(new_n246_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n254_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT72), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n256_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n254_), .B(new_n262_), .C1(new_n255_), .C2(new_n265_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G134gat), .B(G162gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT36), .Z(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n272_), .A2(KEYINPUT36), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n267_), .A2(new_n275_), .A3(new_n268_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(KEYINPUT74), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT37), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n274_), .A2(KEYINPUT74), .A3(KEYINPUT37), .A4(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G57gat), .B(G64gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n283_));
  XOR2_X1   g082(.A(G71gat), .B(G78gat), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n283_), .A2(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G231gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G15gat), .B(G22gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT75), .B(G1gat), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n293_), .A2(G8gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT14), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n292_), .B(new_n297_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n291_), .B(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT17), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n307_), .A2(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n302_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n302_), .A2(KEYINPUT77), .A3(new_n311_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n310_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n281_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n289_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n319_), .B1(new_n233_), .B2(new_n242_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n243_), .A2(KEYINPUT12), .A3(new_n253_), .A4(new_n319_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n251_), .A2(new_n252_), .A3(new_n289_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G230gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT64), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n324_), .A2(KEYINPUT70), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT70), .B1(new_n324_), .B2(new_n327_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n322_), .B(new_n323_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n324_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n326_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G120gat), .B(G148gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT5), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G176gat), .B(G204gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n332_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n336_), .B(KEYINPUT71), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT13), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n330_), .A2(new_n332_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT13), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n337_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n318_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G183gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT25), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G183gat), .ZN(new_n352_));
  INV_X1    g151(.A(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT26), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G190gat), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n350_), .A2(new_n352_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(G169gat), .B2(G176gat), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  INV_X1    g159(.A(G176gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT82), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n362_), .A2(KEYINPUT24), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n367_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n357_), .A2(new_n363_), .A3(KEYINPUT87), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n366_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G218gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G211gat), .ZN(new_n380_));
  INV_X1    g179(.A(G211gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G218gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT21), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G197gat), .B(G204gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G204gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G197gat), .ZN(new_n388_));
  INV_X1    g187(.A(G197gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G204gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(KEYINPUT21), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n384_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n386_), .A2(new_n394_), .B1(new_n383_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n360_), .A2(KEYINPUT22), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT22), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G169gat), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n397_), .A2(new_n399_), .A3(KEYINPUT88), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT88), .B1(new_n397_), .B2(new_n399_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n361_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n349_), .A2(new_n353_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT23), .B1(new_n369_), .B2(new_n371_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n368_), .A2(KEYINPUT23), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n403_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n402_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n378_), .A2(new_n396_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT19), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n385_), .A2(new_n384_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n383_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n393_), .A2(KEYINPUT21), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n415_), .B(new_n416_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n395_), .A2(new_n383_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT86), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n396_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT25), .B(G183gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT26), .B(G190gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n426_), .A2(new_n427_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n370_), .B1(G183gat), .B2(G190gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n368_), .A2(KEYINPUT82), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n367_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n428_), .A2(new_n429_), .B1(new_n432_), .B2(new_n405_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n373_), .B1(new_n364_), .B2(KEYINPUT81), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n372_), .A2(new_n375_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n403_), .ZN(new_n436_));
  AOI21_X1  g235(.A(G176gat), .B1(KEYINPUT83), .B2(KEYINPUT22), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G169gat), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n433_), .A2(new_n434_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n410_), .B(new_n414_), .C1(new_n425_), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n413_), .B1(new_n425_), .B2(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n378_), .A2(new_n409_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n421_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT89), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n446_), .A3(new_n421_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n441_), .B1(new_n448_), .B2(new_n412_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT18), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT90), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  AOI221_X4 g253(.A(KEYINPUT86), .B1(new_n383_), .B2(new_n395_), .C1(new_n386_), .C2(new_n394_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n423_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n436_), .A2(new_n438_), .ZN(new_n458_));
  OAI22_X1  g257(.A1(new_n364_), .A2(KEYINPUT81), .B1(new_n406_), .B2(new_n404_), .ZN(new_n459_));
  OAI22_X1  g258(.A1(new_n428_), .A2(new_n429_), .B1(KEYINPUT24), .B2(new_n362_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n457_), .B2(new_n461_), .ZN(new_n462_));
  AOI211_X1 g261(.A(KEYINPUT89), .B(new_n396_), .C1(new_n378_), .C2(new_n409_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n446_), .B1(new_n443_), .B2(new_n421_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n412_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n440_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n453_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n454_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(KEYINPUT90), .A3(new_n468_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT96), .B(KEYINPUT27), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n477_));
  INV_X1    g276(.A(G141gat), .ZN(new_n478_));
  INV_X1    g277(.A(G148gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT2), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n480_), .A2(new_n483_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n478_), .A2(new_n479_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n481_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT1), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(new_n490_), .A3(new_n475_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n476_), .A2(new_n486_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n493_));
  INV_X1    g292(.A(G127gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(G134gat), .ZN(new_n495_));
  INV_X1    g294(.A(G134gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(G127gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n493_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(G127gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(G134gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT84), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G120gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT84), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT84), .B1(new_n499_), .B2(new_n500_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n492_), .A2(KEYINPUT91), .A3(new_n503_), .A4(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n503_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n486_), .A2(new_n476_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n481_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(G141gat), .A2(G148gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n491_), .A2(new_n513_), .A3(new_n488_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(KEYINPUT91), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n516_), .A3(KEYINPUT4), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G225gat), .A2(G233gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n492_), .A2(KEYINPUT4), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n509_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n508_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n517_), .A2(new_n520_), .A3(KEYINPUT92), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G29gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G57gat), .B(G85gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n523_), .A2(new_n531_), .A3(new_n524_), .A4(new_n525_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G78gat), .B(G106gat), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n510_), .A2(new_n514_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT29), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n421_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(G228gat), .A3(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G228gat), .A2(G233gat), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n422_), .A2(new_n424_), .A3(new_n542_), .A4(new_n539_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n537_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n538_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT28), .B1(new_n538_), .B2(KEYINPUT29), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G22gat), .B(G50gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n547_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n541_), .A2(new_n543_), .A3(new_n537_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n545_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n545_), .B2(new_n554_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n509_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G227gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(G15gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT30), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n439_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n439_), .A2(new_n561_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n557_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G71gat), .B(G99gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G43gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT31), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n439_), .A2(new_n561_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(new_n562_), .A3(new_n509_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n565_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n572_));
  OAI22_X1  g371(.A1(new_n555_), .A2(new_n556_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n568_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n563_), .A2(new_n557_), .A3(new_n564_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n509_), .B1(new_n569_), .B2(new_n562_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n554_), .ZN(new_n578_));
  OAI22_X1  g377(.A1(new_n578_), .A2(new_n544_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n545_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n565_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .A4(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n535_), .B1(new_n573_), .B2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n584_));
  OAI211_X1 g383(.A(new_n410_), .B(new_n584_), .C1(new_n425_), .C2(new_n439_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n412_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n448_), .B2(new_n412_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n468_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n453_), .B(new_n440_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(KEYINPUT27), .A3(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n473_), .A2(new_n583_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(KEYINPUT32), .A3(new_n453_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n453_), .A2(KEYINPUT32), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n449_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n535_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n470_), .A2(new_n471_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n534_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n519_), .A2(new_n509_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n517_), .A2(new_n518_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n508_), .A2(new_n516_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n602_), .B(new_n532_), .C1(new_n603_), .C2(new_n518_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n534_), .B2(new_n599_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n598_), .B1(new_n534_), .B2(new_n599_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n600_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n596_), .B1(new_n597_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n571_), .A2(new_n572_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n555_), .A2(new_n556_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n591_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n247_), .A2(new_n300_), .A3(new_n299_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n246_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT79), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G169gat), .B(G197gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(new_n623_));
  INV_X1    g422(.A(new_n618_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n301_), .A2(new_n246_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(new_n616_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT78), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(KEYINPUT78), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n620_), .B(new_n623_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT80), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n626_), .B(KEYINPUT78), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT80), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n620_), .A4(new_n623_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n620_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n623_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n613_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n348_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT97), .ZN(new_n641_));
  INV_X1    g440(.A(new_n535_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n293_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT38), .ZN(new_n645_));
  INV_X1    g444(.A(G1gat), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n274_), .A2(new_n276_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n613_), .A2(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n338_), .A2(new_n340_), .A3(KEYINPUT13), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n345_), .B1(new_n344_), .B2(new_n337_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n638_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n347_), .A2(KEYINPUT98), .A3(new_n638_), .ZN(new_n655_));
  AND4_X1   g454(.A1(new_n649_), .A2(new_n316_), .A3(new_n654_), .A4(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n646_), .B1(new_n656_), .B2(new_n535_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT99), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n645_), .A2(new_n658_), .ZN(G1324gat));
  INV_X1    g458(.A(G8gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n473_), .A2(new_n590_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n656_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT39), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n641_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g465(.A(new_n559_), .B1(new_n656_), .B2(new_n609_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT41), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n641_), .A2(new_n559_), .A3(new_n609_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1326gat));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n611_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n656_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT42), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n641_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1327gat));
  INV_X1    g475(.A(G29gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT90), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n589_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n449_), .A2(new_n453_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n471_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n607_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n612_), .B1(new_n683_), .B2(new_n595_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n473_), .A2(new_n583_), .A3(new_n590_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n281_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n613_), .A2(new_n688_), .A3(new_n281_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n654_), .A2(new_n317_), .A3(new_n655_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT44), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n694_), .B(new_n691_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n677_), .B1(new_n696_), .B2(new_n535_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n613_), .A2(new_n638_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n699_), .A2(new_n317_), .A3(new_n276_), .A4(new_n274_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n647_), .B2(new_n317_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n698_), .A2(new_n702_), .A3(new_n703_), .A4(new_n347_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n347_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT101), .B1(new_n705_), .B2(new_n639_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(G29gat), .A3(new_n642_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n697_), .A2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(new_n661_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n704_), .A2(new_n706_), .A3(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT45), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT102), .B1(new_n696_), .B2(new_n661_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n613_), .A2(new_n688_), .A3(new_n281_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n688_), .B1(new_n613_), .B2(new_n281_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n692_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n694_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n692_), .B(KEYINPUT44), .C1(new_n715_), .C2(new_n716_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n718_), .A2(KEYINPUT102), .A3(new_n661_), .A4(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT46), .B(new_n713_), .C1(new_n714_), .C2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n713_), .B1(new_n714_), .B2(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT103), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(new_n713_), .C1(new_n714_), .C2(new_n721_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT104), .B(KEYINPUT46), .Z(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AND4_X1   g528(.A1(new_n723_), .A2(new_n725_), .A3(new_n727_), .A4(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n724_), .B2(KEYINPUT103), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n723_), .B1(new_n731_), .B2(new_n727_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n722_), .B1(new_n730_), .B2(new_n732_), .ZN(G1329gat));
  NAND3_X1  g532(.A1(new_n696_), .A2(G43gat), .A3(new_n609_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT106), .B(G43gat), .Z(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n707_), .B2(new_n610_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g537(.A1(new_n696_), .A2(G50gat), .A3(new_n672_), .ZN(new_n739_));
  INV_X1    g538(.A(G50gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n707_), .B2(new_n611_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1331gat));
  INV_X1    g541(.A(new_n638_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n347_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n649_), .A2(new_n316_), .A3(new_n743_), .A4(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT107), .Z(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(G57gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n535_), .A3(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT109), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n347_), .A2(new_n638_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n613_), .A2(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n751_), .A2(new_n317_), .A3(new_n281_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n535_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n749_), .A2(new_n753_), .ZN(G1332gat));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n746_), .B2(new_n661_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT48), .Z(new_n757_));
  NAND3_X1  g556(.A1(new_n752_), .A2(new_n755_), .A3(new_n661_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1333gat));
  INV_X1    g558(.A(G71gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n746_), .B2(new_n609_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT49), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n752_), .A2(new_n760_), .A3(new_n609_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1334gat));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n746_), .B2(new_n672_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT50), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n752_), .A2(new_n765_), .A3(new_n672_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1335gat));
  INV_X1    g568(.A(new_n751_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n702_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n535_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n690_), .A2(new_n317_), .A3(new_n743_), .A4(new_n744_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(KEYINPUT110), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT111), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n535_), .A2(G85gat), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT112), .Z(new_n785_));
  AOI21_X1  g584(.A(new_n773_), .B1(new_n783_), .B2(new_n785_), .ZN(G1336gat));
  NAND2_X1  g585(.A1(new_n661_), .A2(G92gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT113), .Z(new_n788_));
  NAND3_X1  g587(.A1(new_n780_), .A2(new_n782_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G92gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n771_), .B2(new_n710_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(KEYINPUT114), .A3(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n779_), .B2(new_n610_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n772_), .A2(new_n238_), .A3(new_n609_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g599(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n775_), .A2(new_n672_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n803_));
  AND4_X1   g602(.A1(KEYINPUT116), .A2(new_n802_), .A3(G106gat), .A4(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n803_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n222_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n802_), .A2(new_n807_), .B1(KEYINPUT116), .B2(new_n803_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n804_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n772_), .A2(new_n222_), .A3(new_n672_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n801_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n810_), .B(new_n801_), .C1(new_n804_), .C2(new_n808_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  NOR2_X1   g613(.A1(new_n625_), .A2(new_n616_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n619_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n636_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT118), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n636_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n614_), .A2(new_n617_), .A3(new_n816_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n818_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n337_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n330_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n323_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n326_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n330_), .A2(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n343_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n343_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n824_), .B(KEYINPUT58), .C1(new_n831_), .C2(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(new_n281_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n824_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n638_), .A2(new_n337_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n830_), .A2(new_n343_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n343_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n839_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n823_), .B1(new_n340_), .B2(new_n338_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n648_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT57), .B(new_n648_), .C1(new_n844_), .C2(new_n846_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n838_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT54), .B1(new_n348_), .B2(new_n638_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n318_), .A2(new_n853_), .A3(new_n743_), .A4(new_n347_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n851_), .A2(new_n317_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n672_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n661_), .A2(new_n642_), .A3(new_n610_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G113gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n638_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n858_), .A2(new_n861_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n856_), .A2(new_n857_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n743_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n860_), .B1(new_n868_), .B2(new_n859_), .ZN(G1340gat));
  INV_X1    g668(.A(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n347_), .B2(KEYINPUT60), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n870_), .A2(KEYINPUT60), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n856_), .A2(new_n857_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT120), .Z(new_n874_));
  AOI21_X1  g673(.A(new_n347_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n870_), .ZN(G1341gat));
  NAND3_X1  g675(.A1(new_n858_), .A2(new_n494_), .A3(new_n316_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n317_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n494_), .ZN(G1342gat));
  XNOR2_X1  g678(.A(KEYINPUT122), .B(G134gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n281_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n856_), .A2(new_n647_), .A3(new_n857_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(new_n884_), .A3(new_n496_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(new_n496_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n882_), .A2(new_n885_), .A3(new_n886_), .ZN(G1343gat));
  INV_X1    g686(.A(new_n573_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n661_), .A2(new_n642_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n834_), .A2(new_n837_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n316_), .B1(new_n890_), .B2(new_n850_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n852_), .A2(new_n854_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n888_), .B(new_n889_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT123), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n851_), .A2(new_n317_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n892_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n888_), .A4(new_n889_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n638_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n744_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n900_), .B2(new_n316_), .ZN(new_n908_));
  AOI211_X1 g707(.A(KEYINPUT124), .B(new_n317_), .C1(new_n895_), .C2(new_n899_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n573_), .B1(new_n896_), .B2(new_n892_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n898_), .B1(new_n911_), .B2(new_n889_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n889_), .ZN(new_n913_));
  NOR4_X1   g712(.A1(new_n855_), .A2(KEYINPUT123), .A3(new_n573_), .A4(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n316_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT124), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n900_), .A2(new_n907_), .A3(new_n316_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n917_), .A3(new_n905_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n918_), .ZN(G1346gat));
  INV_X1    g718(.A(new_n900_), .ZN(new_n920_));
  OR3_X1    g719(.A1(new_n920_), .A2(G162gat), .A3(new_n648_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n281_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G162gat), .B1(new_n920_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n710_), .A2(new_n535_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n610_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n856_), .A2(new_n927_), .ZN(new_n928_));
  AOI211_X1 g727(.A(KEYINPUT62), .B(new_n360_), .C1(new_n928_), .C2(new_n638_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n638_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(G169gat), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n928_), .B(new_n638_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n929_), .B1(new_n932_), .B2(new_n933_), .ZN(G1348gat));
  NAND2_X1  g733(.A1(new_n928_), .A2(new_n744_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g735(.A(new_n426_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n928_), .A2(new_n937_), .A3(new_n316_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n938_), .A2(KEYINPUT125), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(KEYINPUT125), .ZN(new_n940_));
  AOI21_X1  g739(.A(G183gat), .B1(new_n928_), .B2(new_n316_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n941_), .ZN(G1350gat));
  INV_X1    g741(.A(new_n928_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G190gat), .B1(new_n943_), .B2(new_n922_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n928_), .A2(new_n647_), .A3(new_n427_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1351gat));
  NOR3_X1   g745(.A1(new_n855_), .A2(new_n573_), .A3(new_n926_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n638_), .ZN(new_n948_));
  XOR2_X1   g747(.A(KEYINPUT126), .B(G197gat), .Z(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1352gat));
  NAND2_X1  g749(.A1(new_n947_), .A2(new_n744_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  NAND2_X1  g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n947_), .A2(new_n316_), .A3(new_n953_), .A4(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n947_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n317_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n955_), .B1(new_n959_), .B2(new_n953_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n957_), .B1(new_n960_), .B2(KEYINPUT127), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n958_), .B2(new_n922_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n947_), .A2(new_n379_), .A3(new_n647_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1355gat));
endmodule


