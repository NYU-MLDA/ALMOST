//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n847_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_;
  NOR2_X1   g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT65), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  AND2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n209_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n205_), .A2(KEYINPUT65), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n204_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G85gat), .B(G92gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT68), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT69), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(new_n223_), .A3(new_n210_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n224_), .A3(new_n204_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n217_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT8), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n225_), .B2(new_n217_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n219_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(G92gat), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT9), .ZN(new_n233_));
  INV_X1    g032(.A(new_n216_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(KEYINPUT9), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT10), .B(G99gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(G106gat), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n214_), .A2(new_n210_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT71), .Z(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(KEYINPUT11), .B2(new_n241_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n243_), .B(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n230_), .A2(new_n240_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT72), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n230_), .A2(new_n240_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n246_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n230_), .A2(KEYINPUT72), .A3(new_n240_), .A4(new_n246_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT64), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n225_), .A2(new_n217_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT70), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT8), .A3(new_n227_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n239_), .B1(new_n260_), .B2(new_n219_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n256_), .B1(new_n261_), .B2(new_n246_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n264_));
  AOI211_X1 g063(.A(KEYINPUT12), .B(new_n246_), .C1(new_n230_), .C2(new_n240_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n262_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G120gat), .B(G148gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G176gat), .B(G204gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n257_), .A2(new_n266_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT74), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n257_), .A2(new_n266_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n271_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(KEYINPUT74), .A3(new_n273_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n276_), .A2(new_n279_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G29gat), .B(G36gat), .Z(new_n289_));
  XOR2_X1   g088(.A(G43gat), .B(G50gat), .Z(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT15), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n292_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G229gat), .A2(G233gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n291_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(new_n300_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n291_), .B(new_n299_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n301_), .A2(new_n305_), .B1(new_n306_), .B2(new_n303_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G113gat), .B(G141gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(G169gat), .B(G197gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n307_), .A2(new_n310_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n288_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT89), .B(G197gat), .Z(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(G204gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G211gat), .B(G218gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT89), .B(G197gat), .ZN(new_n323_));
  INV_X1    g122(.A(G204gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT90), .B1(new_n325_), .B2(new_n317_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n321_), .A2(KEYINPUT21), .A3(new_n322_), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n324_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(G197gat), .B2(G204gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n322_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(KEYINPUT21), .B2(new_n319_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n341_));
  OAI22_X1  g140(.A1(new_n339_), .A2(new_n340_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n336_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n340_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n337_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT25), .B(G183gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n349_), .A2(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G176gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT24), .B1(new_n335_), .B2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(new_n352_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n345_), .B1(new_n348_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n316_), .B1(new_n333_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n327_), .A2(new_n332_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n352_), .B1(new_n355_), .B2(KEYINPUT94), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(KEYINPUT94), .B2(new_n355_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(new_n342_), .A3(new_n353_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT95), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n362_), .A2(new_n342_), .A3(KEYINPUT95), .A4(new_n353_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT96), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n348_), .A2(new_n368_), .A3(new_n344_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n339_), .A2(new_n340_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT96), .B1(new_n370_), .B2(new_n343_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n336_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n360_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT19), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n359_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n327_), .A2(new_n332_), .A3(new_n363_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n378_), .B2(new_n372_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT100), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n357_), .A2(new_n348_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n342_), .A2(new_n344_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(new_n336_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n360_), .ZN(new_n385_));
  OAI211_X1 g184(.A(KEYINPUT100), .B(KEYINPUT20), .C1(new_n378_), .C2(new_n372_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n381_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n377_), .B1(new_n387_), .B2(new_n375_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G8gat), .B(G36gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n369_), .A2(new_n371_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n336_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(new_n333_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n376_), .A2(KEYINPUT20), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n384_), .B2(new_n360_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT20), .B1(new_n384_), .B2(new_n360_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n398_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n360_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n394_), .B(new_n402_), .C1(new_n405_), .C2(new_n376_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT27), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n395_), .A2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n399_), .A2(new_n401_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n376_), .B1(new_n359_), .B2(new_n373_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n393_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n406_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT27), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT103), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT103), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n408_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G141gat), .A2(G148gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT3), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT2), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424_));
  OR2_X1    g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT87), .B1(new_n424_), .B2(KEYINPUT1), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(G155gat), .A4(G162gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(KEYINPUT1), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n427_), .A2(new_n430_), .A3(new_n425_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n433_));
  XOR2_X1   g232(.A(G141gat), .B(G148gat), .Z(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n433_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n426_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n440_));
  OAI21_X1  g239(.A(new_n360_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n442_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n438_), .A2(KEYINPUT29), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(KEYINPUT91), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT91), .B1(new_n446_), .B2(new_n447_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n443_), .B(new_n445_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n443_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n444_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n438_), .A2(KEYINPUT29), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G22gat), .B(G50gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT28), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n455_), .B(new_n457_), .ZN(new_n458_));
  AND4_X1   g257(.A1(new_n451_), .A2(new_n452_), .A3(new_n454_), .A4(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n452_), .A2(new_n458_), .B1(new_n454_), .B2(new_n451_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G127gat), .B(G134gat), .Z(new_n462_));
  XOR2_X1   g261(.A(G113gat), .B(G120gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT83), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT84), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G127gat), .B(G134gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G113gat), .B(G120gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n464_), .A2(KEYINPUT83), .A3(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n466_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n438_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n464_), .A2(new_n469_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT98), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n439_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n475_), .A2(new_n478_), .A3(KEYINPUT4), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT4), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n482_), .B(new_n438_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n479_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n480_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G1gat), .B(G29gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G85gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n491_), .B(new_n480_), .C1(new_n481_), .C2(new_n485_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT102), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(KEYINPUT102), .A3(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n358_), .B(KEYINPUT30), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT82), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n384_), .B(KEYINPUT30), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT82), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G71gat), .B(G99gat), .ZN(new_n507_));
  INV_X1    g306(.A(G43gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(G15gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n509_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n473_), .A2(new_n474_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n516_), .A2(KEYINPUT85), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(KEYINPUT85), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT31), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n505_), .A2(new_n513_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT31), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n515_), .A2(new_n519_), .A3(new_n520_), .A4(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n520_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n513_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n519_), .ZN(new_n526_));
  OAI22_X1  g325(.A1(new_n524_), .A2(new_n525_), .B1(new_n526_), .B2(new_n521_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n418_), .A2(new_n461_), .A3(new_n500_), .A4(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n461_), .A2(new_n499_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n394_), .A2(KEYINPUT32), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n409_), .A2(new_n410_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT101), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n388_), .B2(new_n531_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n386_), .A2(new_n385_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n376_), .B1(new_n537_), .B2(new_n381_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT101), .B(new_n532_), .C1(new_n538_), .C2(new_n377_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n494_), .B(KEYINPUT33), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n475_), .A2(new_n478_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n483_), .A2(new_n479_), .ZN(new_n543_));
  OAI221_X1 g342(.A(new_n492_), .B1(new_n479_), .B2(new_n542_), .C1(new_n481_), .C2(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n544_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n530_), .A2(new_n418_), .B1(new_n547_), .B2(new_n461_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT86), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n528_), .B(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n529_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n250_), .A2(new_n292_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n250_), .A2(new_n304_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n558_), .A2(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n555_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n250_), .A2(new_n292_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n261_), .A2(new_n291_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT77), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n562_), .A2(new_n564_), .A3(KEYINPUT76), .A4(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n563_), .A2(new_n555_), .B1(new_n568_), .B2(KEYINPUT77), .ZN(new_n576_));
  INV_X1    g375(.A(new_n574_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n576_), .A2(KEYINPUT76), .A3(new_n577_), .A4(new_n562_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n562_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n575_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT37), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n299_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n246_), .B(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G127gat), .B(G155gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n586_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n593_), .B2(new_n586_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT79), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n575_), .A2(new_n581_), .A3(new_n598_), .A4(new_n578_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n583_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n315_), .A2(new_n552_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n294_), .A3(new_n499_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n315_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n582_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n551_), .A2(new_n597_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n500_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n603_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n609_), .A3(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n418_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n601_), .A2(new_n295_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  INV_X1    g413(.A(new_n608_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n612_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n616_), .B2(G8gat), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT39), .B(new_n295_), .C1(new_n615_), .C2(new_n612_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n613_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(G1325gat));
  INV_X1    g420(.A(new_n550_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G15gat), .B1(new_n608_), .B2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT41), .Z(new_n624_));
  NAND3_X1  g423(.A1(new_n601_), .A2(new_n511_), .A3(new_n550_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1326gat));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n461_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n601_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n615_), .B2(new_n628_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n597_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n551_), .A2(new_n635_), .A3(new_n582_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n315_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G29gat), .A3(new_n500_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n284_), .A2(new_n287_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(new_n313_), .A3(new_n597_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n583_), .A2(new_n599_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT43), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n551_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n551_), .B2(new_n642_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT44), .B(new_n641_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n499_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n639_), .B1(new_n652_), .B2(G29gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT105), .ZN(G1328gat));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  INV_X1    g454(.A(new_n636_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n418_), .A2(G36gat), .ZN(new_n657_));
  AND4_X1   g456(.A1(new_n655_), .A2(new_n605_), .A3(new_n656_), .A4(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n637_), .B2(new_n657_), .ZN(new_n659_));
  OAI22_X1  g458(.A1(new_n658_), .A2(new_n659_), .B1(KEYINPUT107), .B2(KEYINPUT46), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n650_), .A2(new_n612_), .A3(new_n651_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(G36gat), .B2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT107), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n662_), .B(new_n664_), .ZN(G1329gat));
  NAND4_X1  g464(.A1(new_n650_), .A2(G43gat), .A3(new_n528_), .A4(new_n651_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n508_), .B1(new_n638_), .B2(new_n622_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g468(.A1(new_n638_), .A2(G50gat), .A3(new_n461_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n650_), .A2(KEYINPUT108), .A3(new_n628_), .A4(new_n651_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(G50gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n650_), .A2(new_n628_), .A3(new_n651_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT109), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  AND4_X1   g475(.A1(KEYINPUT109), .A2(new_n675_), .A3(G50gat), .A4(new_n671_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n670_), .B1(new_n676_), .B2(new_n677_), .ZN(G1331gat));
  NOR2_X1   g477(.A1(new_n288_), .A2(new_n314_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n607_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n500_), .ZN(new_n682_));
  NOR4_X1   g481(.A1(new_n552_), .A2(new_n288_), .A3(new_n314_), .A4(new_n600_), .ZN(new_n683_));
  INV_X1    g482(.A(G57gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n499_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1332gat));
  INV_X1    g485(.A(G64gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n680_), .B2(new_n612_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n683_), .A2(new_n687_), .A3(new_n612_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1333gat));
  INV_X1    g491(.A(G71gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n683_), .A2(new_n693_), .A3(new_n550_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT49), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n680_), .A2(new_n550_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(G71gat), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT49), .B(new_n693_), .C1(new_n680_), .C2(new_n550_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT111), .ZN(G1334gat));
  INV_X1    g499(.A(G78gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n680_), .B2(new_n628_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n683_), .A2(new_n701_), .A3(new_n628_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1335gat));
  NOR3_X1   g505(.A1(new_n288_), .A2(new_n314_), .A3(new_n597_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n231_), .B1(new_n709_), .B2(new_n499_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n656_), .A2(new_n679_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT113), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n499_), .A2(new_n231_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT114), .ZN(G1336gat));
  OAI21_X1  g515(.A(G92gat), .B1(new_n708_), .B2(new_n418_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n612_), .A2(new_n232_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n713_), .B2(new_n718_), .ZN(G1337gat));
  OAI21_X1  g518(.A(G99gat), .B1(new_n708_), .B2(new_n622_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n528_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n236_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n713_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g524(.A1(new_n709_), .A2(new_n628_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(G106gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G106gat), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n461_), .A2(G106gat), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n728_), .A2(new_n729_), .B1(new_n713_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT53), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n733_));
  OAI221_X1 g532(.A(new_n733_), .B1(new_n713_), .B2(new_n730_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1339gat));
  OAI211_X1 g534(.A(new_n301_), .B(new_n303_), .C1(new_n299_), .C2(new_n291_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n310_), .B1(new_n306_), .B2(new_n302_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n311_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n279_), .A2(new_n276_), .A3(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n314_), .A2(new_n273_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n264_), .A2(new_n265_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n249_), .A2(new_n253_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n256_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n266_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT55), .B(new_n262_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n741_), .B1(new_n748_), .B2(new_n271_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n740_), .B1(new_n749_), .B2(KEYINPUT56), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n741_), .B(new_n751_), .C1(new_n748_), .C2(new_n271_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n739_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n606_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT57), .A3(new_n606_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n748_), .A2(new_n271_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n751_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n273_), .A2(new_n738_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n748_), .A2(KEYINPUT56), .A3(new_n271_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT116), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT56), .B1(new_n748_), .B2(new_n271_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n760_), .B(new_n761_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n758_), .A2(new_n751_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(KEYINPUT116), .A3(new_n762_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n766_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n760_), .A4(new_n761_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(new_n642_), .A3(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n756_), .A2(new_n757_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n635_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n284_), .A2(new_n313_), .A3(new_n287_), .ZN(new_n775_));
  OR3_X1    g574(.A1(new_n775_), .A2(new_n600_), .A3(KEYINPUT54), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT54), .B1(new_n775_), .B2(new_n600_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n612_), .A2(new_n721_), .A3(new_n628_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n499_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G113gat), .B1(new_n784_), .B2(new_n314_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT59), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n773_), .A2(new_n635_), .B1(new_n777_), .B2(new_n776_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n781_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n765_), .A2(new_n766_), .B1(new_n599_), .B2(new_n583_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n771_), .A2(new_n789_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n597_), .B1(new_n790_), .B2(new_n757_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n776_), .A2(new_n777_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT59), .B(new_n782_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n788_), .A2(new_n793_), .A3(KEYINPUT118), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT118), .B1(new_n788_), .B2(new_n793_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n314_), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(KEYINPUT119), .B2(G113gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n785_), .B1(new_n796_), .B2(new_n798_), .ZN(G1340gat));
  NAND2_X1  g598(.A1(new_n788_), .A2(new_n793_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT120), .B(G120gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n640_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT60), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n288_), .B1(new_n784_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n784_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n800_), .A2(new_n805_), .B1(new_n806_), .B2(new_n801_), .ZN(G1341gat));
  AOI21_X1  g606(.A(G127gat), .B1(new_n784_), .B2(new_n597_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n597_), .A2(G127gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n796_), .B2(new_n809_), .ZN(G1342gat));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n787_), .A2(new_n606_), .A3(new_n781_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(G134gat), .ZN(new_n813_));
  INV_X1    g612(.A(G134gat), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT121), .B(new_n814_), .C1(new_n783_), .C2(new_n606_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n642_), .ZN(new_n817_));
  XOR2_X1   g616(.A(KEYINPUT122), .B(G134gat), .Z(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n816_), .B1(new_n796_), .B2(new_n819_), .ZN(G1343gat));
  NOR4_X1   g619(.A1(new_n550_), .A2(new_n612_), .A3(new_n461_), .A4(new_n500_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT123), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n779_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n314_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n640_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g627(.A1(new_n823_), .A2(new_n635_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT61), .B(G155gat), .Z(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  OR3_X1    g630(.A1(new_n823_), .A2(G162gat), .A3(new_n606_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G162gat), .B1(new_n823_), .B2(new_n817_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1347gat));
  INV_X1    g633(.A(KEYINPUT22), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n622_), .A2(new_n628_), .A3(new_n499_), .A4(new_n418_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n779_), .A2(new_n835_), .A3(new_n314_), .A4(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT62), .A3(new_n335_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(KEYINPUT62), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n779_), .A2(new_n314_), .A3(new_n836_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G169gat), .B1(new_n840_), .B2(KEYINPUT62), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(G1348gat));
  NAND2_X1  g642(.A1(new_n779_), .A2(new_n836_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n288_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n354_), .ZN(G1349gat));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n635_), .ZN(new_n847_));
  MUX2_X1   g646(.A(G183gat), .B(new_n349_), .S(new_n847_), .Z(G1350gat));
  OAI21_X1  g647(.A(G190gat), .B1(new_n844_), .B2(new_n817_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n582_), .A2(new_n350_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n844_), .B2(new_n850_), .ZN(G1351gat));
  XNOR2_X1  g650(.A(KEYINPUT124), .B(G197gat), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(G197gat), .ZN(new_n854_));
  NOR4_X1   g653(.A1(new_n550_), .A2(new_n461_), .A3(new_n499_), .A4(new_n418_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n779_), .A2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n313_), .ZN(new_n857_));
  MUX2_X1   g656(.A(new_n852_), .B(new_n854_), .S(new_n857_), .Z(G1352gat));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n288_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(KEYINPUT125), .B2(new_n324_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT125), .B(G204gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n859_), .B2(new_n861_), .ZN(G1353gat));
  INV_X1    g661(.A(new_n856_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n635_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT126), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n865_), .B(new_n867_), .ZN(G1354gat));
  OR3_X1    g667(.A1(new_n856_), .A2(G218gat), .A3(new_n606_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G218gat), .B1(new_n856_), .B2(new_n817_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1355gat));
endmodule


