//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G232gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT34), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT35), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n210_), .A2(KEYINPUT75), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT10), .B(G99gat), .Z(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n221_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT9), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(G85gat), .B2(G92gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT66), .B(new_n220_), .C1(new_n228_), .C2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT67), .B1(G85gat), .B2(G92gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n234_), .B1(new_n237_), .B2(new_n217_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT8), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n231_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n220_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n232_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G43gat), .B(G50gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(G29gat), .B(G36gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n207_), .A2(KEYINPUT35), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(KEYINPUT69), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n247_), .B(KEYINPUT15), .Z(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n232_), .A2(new_n239_), .A3(new_n243_), .A4(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  AOI211_X1 g054(.A(new_n213_), .B(new_n214_), .C1(new_n250_), .C2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n250_), .A2(new_n255_), .A3(KEYINPUT75), .A4(new_n210_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n205_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT76), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT76), .B(new_n205_), .C1(new_n256_), .C2(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n214_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n213_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n204_), .B(KEYINPUT36), .Z(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n257_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT37), .B1(new_n263_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT37), .ZN(new_n270_));
  INV_X1    g069(.A(new_n268_), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n270_), .B(new_n271_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT77), .B(G15gat), .ZN(new_n274_));
  INV_X1    g073(.A(G22gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G1gat), .ZN(new_n277_));
  INV_X1    g076(.A(G8gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT14), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n281_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(G231gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G57gat), .B(G64gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT11), .ZN(new_n288_));
  XOR2_X1   g087(.A(G71gat), .B(G78gat), .Z(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n288_), .A2(new_n289_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n287_), .A2(KEYINPUT11), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n286_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G127gat), .B(G155gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT16), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G183gat), .B(G211gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT17), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n298_), .B(new_n303_), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n296_), .A2(KEYINPUT17), .A3(new_n302_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n273_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT79), .Z(new_n308_));
  NAND4_X1  g107(.A1(new_n232_), .A2(new_n239_), .A3(new_n243_), .A4(new_n295_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT68), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT68), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n244_), .A2(new_n294_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n294_), .A2(KEYINPUT12), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n251_), .A2(new_n254_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT12), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n312_), .A2(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n309_), .A2(KEYINPUT70), .A3(new_n314_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT70), .B1(new_n309_), .B2(new_n314_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n319_), .B(new_n321_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT72), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G120gat), .B(G148gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G176gat), .B(G204gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NAND3_X1  g129(.A1(new_n316_), .A2(new_n324_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT73), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n316_), .B2(new_n324_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT13), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT13), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(KEYINPUT74), .A3(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n308_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT22), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT22), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G169gat), .ZN(new_n349_));
  INV_X1    g148(.A(G176gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356_));
  INV_X1    g155(.A(G183gat), .ZN(new_n357_));
  INV_X1    g156(.A(G190gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n359_), .B(new_n360_), .C1(G183gat), .C2(G190gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n351_), .A2(KEYINPUT82), .A3(new_n352_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(KEYINPUT24), .A3(new_n366_), .A4(new_n352_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n359_), .A2(new_n360_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT25), .B(G183gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT24), .ZN(new_n372_));
  INV_X1    g171(.A(new_n366_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n364_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n367_), .A2(new_n368_), .A3(new_n371_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n363_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(G15gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G71gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(G99gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n377_), .B(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G127gat), .B(G134gat), .Z(new_n384_));
  XOR2_X1   g183(.A(G113gat), .B(G120gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n383_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT83), .B(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT31), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n390_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G141gat), .ZN(new_n394_));
  INV_X1    g193(.A(G148gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(KEYINPUT84), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(G141gat), .B2(G148gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n399_), .A2(new_n402_), .A3(new_n405_), .A4(KEYINPUT85), .ZN(new_n409_));
  NOR2_X1   g208(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n411_));
  OAI22_X1  g210(.A1(KEYINPUT86), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT2), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n401_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G155gat), .B(G162gat), .Z(new_n417_));
  AOI22_X1  g216(.A1(new_n408_), .A2(new_n409_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n420_), .B(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G22gat), .B(G50gat), .Z(new_n424_));
  AND2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n423_), .A2(new_n424_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT88), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT90), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n416_), .A2(new_n417_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n400_), .A2(new_n401_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n398_), .B2(new_n396_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT85), .B1(new_n433_), .B2(new_n405_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n409_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n431_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT29), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT21), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  AND2_X1   g238(.A1(G197gat), .A2(G204gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G197gat), .A2(G204gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G211gat), .B(G218gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G218gat), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n445_), .A2(G211gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(G211gat), .ZN(new_n447_));
  OAI22_X1  g246(.A1(new_n446_), .A2(new_n447_), .B1(new_n441_), .B2(new_n440_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n438_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT21), .B1(new_n442_), .B2(new_n443_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n430_), .B1(new_n437_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT90), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n429_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n451_), .B(new_n454_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n452_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n430_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n408_), .A2(new_n409_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n419_), .B1(new_n460_), .B2(new_n431_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n451_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n463_), .A2(KEYINPUT91), .A3(new_n455_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT91), .B1(new_n463_), .B2(new_n455_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n457_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n458_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n457_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n463_), .A2(KEYINPUT91), .A3(new_n455_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT92), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n427_), .B1(new_n468_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n458_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n469_), .B1(new_n463_), .B2(new_n455_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT93), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n425_), .A2(new_n426_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n476_), .B1(new_n473_), .B2(KEYINPUT92), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n466_), .A2(new_n467_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n477_), .A2(new_n478_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n376_), .A2(new_n451_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n352_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT22), .B(G169gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(new_n350_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n353_), .A2(KEYINPUT94), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n361_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n372_), .A2(new_n346_), .A3(new_n350_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n367_), .A2(new_n371_), .A3(new_n368_), .A4(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n495_), .B(new_n497_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT19), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AND4_X1   g300(.A1(KEYINPUT20), .A2(new_n488_), .A3(new_n498_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT20), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n361_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n353_), .A2(KEYINPUT94), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n497_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n503_), .B1(new_n506_), .B2(new_n451_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n363_), .B(new_n375_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n501_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G8gat), .B(G36gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n502_), .A2(new_n509_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n506_), .A2(new_n451_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n508_), .A3(KEYINPUT20), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n500_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n488_), .A2(new_n498_), .A3(KEYINPUT20), .A4(new_n501_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n516_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n515_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT27), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT99), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n488_), .A2(new_n498_), .A3(KEYINPUT20), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n500_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n507_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT99), .B1(new_n525_), .B2(new_n500_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n514_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n515_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT27), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G225gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT96), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n436_), .A2(new_n537_), .A3(new_n387_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n436_), .A2(new_n387_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n418_), .A2(new_n386_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n536_), .B(new_n538_), .C1(new_n541_), .C2(new_n537_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n536_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G1gat), .B(G29gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G57gat), .B(G85gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n542_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n480_), .A2(new_n487_), .A3(new_n534_), .A4(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n521_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n543_), .B(new_n538_), .C1(new_n541_), .C2(new_n537_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n558_), .B(new_n551_), .C1(new_n543_), .C2(new_n541_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n531_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT98), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n542_), .A2(new_n544_), .A3(KEYINPUT33), .A4(new_n550_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .A4(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n522_), .A2(new_n563_), .A3(new_n564_), .A4(new_n559_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n519_), .A2(new_n520_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n516_), .A2(KEYINPUT32), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n552_), .A2(new_n553_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT32), .B(new_n516_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n566_), .A2(KEYINPUT98), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n480_), .A2(new_n487_), .B1(new_n565_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n556_), .B1(new_n573_), .B2(KEYINPUT100), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575_));
  AOI221_X4 g374(.A(new_n575_), .B1(new_n572_), .B2(new_n565_), .C1(new_n480_), .C2(new_n487_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n393_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n475_), .A2(KEYINPUT93), .A3(new_n479_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n485_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n393_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(new_n555_), .A4(new_n534_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT101), .B(new_n393_), .C1(new_n574_), .C2(new_n576_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT80), .B1(new_n284_), .B2(new_n247_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT80), .ZN(new_n589_));
  INV_X1    g388(.A(new_n247_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n282_), .A2(new_n589_), .A3(new_n283_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n284_), .A2(new_n247_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n588_), .A2(new_n591_), .B1(new_n284_), .B2(new_n252_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n596_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n596_), .B(new_n603_), .C1(new_n594_), .C2(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n587_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n345_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n607_), .A2(G1gat), .A3(new_n555_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT38), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT38), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n342_), .A2(new_n605_), .A3(new_n343_), .A4(new_n306_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT102), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n263_), .A2(new_n268_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT103), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n587_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n555_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n609_), .A2(new_n610_), .A3(new_n618_), .ZN(G1324gat));
  INV_X1    g418(.A(new_n607_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n278_), .A3(new_n533_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n612_), .A2(new_n616_), .A3(new_n533_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n621_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g427(.A(G15gat), .B1(new_n617_), .B2(new_n393_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT105), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n620_), .A2(new_n379_), .A3(new_n584_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(G1326gat));
  NAND3_X1  g434(.A1(new_n620_), .A2(new_n275_), .A3(new_n582_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n612_), .A2(new_n616_), .A3(new_n582_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT42), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(G22gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n637_), .B2(G22gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n636_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT106), .ZN(G1327gat));
  INV_X1    g442(.A(new_n344_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n613_), .A2(new_n306_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n587_), .A2(new_n644_), .A3(new_n605_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n554_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n605_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n344_), .A2(new_n649_), .A3(new_n306_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  INV_X1    g450(.A(new_n273_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n586_), .A2(new_n585_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n572_), .A2(new_n565_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n575_), .B1(new_n582_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n573_), .A2(KEYINPUT100), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n556_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT101), .B1(new_n657_), .B2(new_n393_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n651_), .B(new_n652_), .C1(new_n653_), .C2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n651_), .B1(new_n587_), .B2(new_n652_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n650_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT44), .B(new_n650_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n554_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n648_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n533_), .A3(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G36gat), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n646_), .A2(G36gat), .A3(new_n534_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT45), .Z(new_n672_));
  OR2_X1    g471(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1329gat));
  AOI21_X1  g475(.A(G43gat), .B1(new_n647_), .B2(new_n584_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n584_), .A2(G43gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n666_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT47), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1330gat));
  OR3_X1    g480(.A1(new_n646_), .A2(G50gat), .A3(new_n583_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n664_), .A2(new_n683_), .A3(new_n582_), .A4(new_n665_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(G50gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n664_), .A2(new_n582_), .A3(new_n665_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT108), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT109), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  AND4_X1   g487(.A1(KEYINPUT109), .A2(new_n687_), .A3(G50gat), .A4(new_n684_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n682_), .B1(new_n688_), .B2(new_n689_), .ZN(G1331gat));
  NAND2_X1  g489(.A1(new_n306_), .A2(new_n649_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n616_), .A2(new_n344_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G57gat), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n555_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT110), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n308_), .A2(new_n644_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n587_), .A2(new_n649_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n694_), .B1(new_n700_), .B2(new_n555_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n696_), .A2(KEYINPUT110), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n697_), .A2(new_n701_), .A3(new_n702_), .ZN(G1332gat));
  OAI21_X1  g502(.A(G64gat), .B1(new_n693_), .B2(new_n534_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT48), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n534_), .A2(G64gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n700_), .B2(new_n706_), .ZN(G1333gat));
  OAI21_X1  g506(.A(G71gat), .B1(new_n693_), .B2(new_n393_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT49), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n393_), .A2(G71gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n700_), .B2(new_n710_), .ZN(G1334gat));
  OAI21_X1  g510(.A(G78gat), .B1(new_n693_), .B2(new_n583_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n583_), .A2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n700_), .B2(new_n714_), .ZN(G1335gat));
  AND2_X1   g514(.A1(new_n344_), .A2(new_n645_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n699_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n554_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT111), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n660_), .A2(new_n661_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n306_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n344_), .A2(new_n649_), .A3(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT112), .Z(new_n724_));
  AND2_X1   g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n554_), .A2(G85gat), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT113), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n720_), .B1(new_n725_), .B2(new_n727_), .ZN(G1336gat));
  INV_X1    g527(.A(G92gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n718_), .A2(new_n729_), .A3(new_n533_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n725_), .A2(new_n533_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n729_), .ZN(G1337gat));
  NAND2_X1  g531(.A1(new_n584_), .A2(new_n219_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734_));
  OAI22_X1  g533(.A1(new_n717_), .A2(new_n733_), .B1(KEYINPUT114), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n725_), .A2(new_n584_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G99gat), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n734_), .A2(KEYINPUT114), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n718_), .A2(new_n218_), .A3(new_n582_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n721_), .A2(new_n724_), .A3(new_n582_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G106gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT53), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(new_n740_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1339gat));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(KEYINPUT54), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n340_), .A2(new_n692_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n652_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n751_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n340_), .A2(new_n273_), .A3(new_n692_), .A4(new_n754_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n753_), .A2(new_n755_), .B1(new_n750_), .B2(KEYINPUT54), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n592_), .A2(new_n595_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n601_), .B1(new_n757_), .B2(new_n593_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n597_), .A2(new_n594_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n598_), .A2(new_n601_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n331_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n330_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n319_), .A2(new_n309_), .A3(new_n321_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n315_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(KEYINPUT118), .A3(new_n315_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n766_), .B(new_n767_), .C1(new_n768_), .C2(new_n324_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n324_), .A2(KEYINPUT117), .A3(new_n768_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT117), .B1(new_n324_), .B2(new_n768_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n762_), .B1(new_n769_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n324_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n776_), .A2(KEYINPUT55), .B1(new_n764_), .B2(new_n765_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n767_), .C1(new_n771_), .C2(new_n770_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n762_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n761_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n781_));
  AOI21_X1  g580(.A(new_n273_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT120), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n773_), .A2(new_n774_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n762_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(KEYINPUT58), .A4(new_n761_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(new_n784_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n605_), .A2(new_n331_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n605_), .A2(KEYINPUT116), .A3(new_n331_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n336_), .A2(new_n760_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n613_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT57), .B(new_n613_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n790_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n756_), .B1(new_n802_), .B2(new_n722_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n393_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n582_), .A2(new_n555_), .A3(new_n533_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n605_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n649_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n813_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n644_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n807_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n644_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n815_), .ZN(G1341gat));
  INV_X1    g618(.A(G127gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n807_), .A2(new_n820_), .A3(new_n306_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n722_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n820_), .ZN(G1342gat));
  AOI21_X1  g622(.A(G134gat), .B1(new_n807_), .B2(new_n614_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n810_), .A2(new_n812_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT121), .B(G134gat), .Z(new_n826_));
  NOR2_X1   g625(.A1(new_n273_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(G1343gat));
  NAND2_X1  g627(.A1(new_n802_), .A2(new_n722_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n756_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n583_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AND4_X1   g630(.A1(new_n393_), .A2(new_n831_), .A3(new_n554_), .A4(new_n534_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n605_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n344_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n306_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1346gat));
  INV_X1    g638(.A(G162gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n832_), .A2(new_n840_), .A3(new_n614_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n832_), .A2(new_n652_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n840_), .ZN(G1347gat));
  NOR2_X1   g642(.A1(new_n534_), .A2(new_n554_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n582_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n804_), .A2(new_n605_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT122), .B1(new_n847_), .B2(G169gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n804_), .A2(new_n846_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n605_), .A3(new_n490_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n849_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(new_n855_), .A3(new_n856_), .ZN(G1348gat));
  NOR2_X1   g656(.A1(new_n853_), .A2(new_n644_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT123), .B(G176gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1349gat));
  NAND2_X1  g659(.A1(new_n854_), .A2(new_n306_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(G183gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n369_), .B1(KEYINPUT124), .B2(G183gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n861_), .B2(new_n864_), .ZN(G1350gat));
  OAI21_X1  g664(.A(G190gat), .B1(new_n853_), .B2(new_n273_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n614_), .A2(new_n370_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n853_), .B2(new_n867_), .ZN(G1351gat));
  NOR2_X1   g667(.A1(new_n845_), .A2(new_n584_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n800_), .A2(new_n801_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n306_), .B1(new_n870_), .B2(new_n790_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n582_), .B(new_n869_), .C1(new_n871_), .C2(new_n756_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT125), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n831_), .A2(new_n874_), .A3(new_n869_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n605_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g677(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT126), .B(G204gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n344_), .ZN(new_n881_));
  MUX2_X1   g680(.A(new_n879_), .B(new_n880_), .S(new_n881_), .Z(G1353gat));
  OR2_X1    g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  AND4_X1   g683(.A1(new_n306_), .A2(new_n876_), .A3(new_n883_), .A4(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n876_), .B2(new_n306_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1354gat));
  AOI21_X1  g686(.A(new_n874_), .B1(new_n831_), .B2(new_n869_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n869_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n803_), .A2(KEYINPUT125), .A3(new_n583_), .A4(new_n889_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n445_), .B(new_n614_), .C1(new_n888_), .C2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT127), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n273_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n892_), .C1(new_n893_), .C2(new_n445_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n652_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G218gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n892_), .B1(new_n897_), .B2(new_n891_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1355gat));
endmodule


