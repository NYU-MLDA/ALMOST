//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT64), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G57gat), .B(G64gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n207_));
  XOR2_X1   g006(.A(G71gat), .B(G78gat), .Z(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(KEYINPUT65), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(KEYINPUT65), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(G99gat), .A4(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(KEYINPUT66), .A3(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n238_));
  INV_X1    g037(.A(G99gat), .ZN(new_n239_));
  INV_X1    g038(.A(G106gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n219_), .B1(new_n233_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n243_), .A2(new_n246_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n237_), .A2(new_n242_), .A3(KEYINPUT68), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n216_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n218_), .B1(new_n249_), .B2(KEYINPUT69), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n241_), .B1(new_n251_), .B2(new_n238_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n234_), .A2(new_n236_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n246_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n248_), .A3(new_n229_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n217_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n245_), .B1(new_n250_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n216_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT10), .B(G99gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(G106gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n261_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n233_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n209_), .B(new_n211_), .C1(new_n259_), .C2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n233_), .A2(new_n244_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n219_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n255_), .A2(KEYINPUT69), .A3(new_n217_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT8), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n255_), .B2(new_n217_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n211_), .A2(new_n209_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n266_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n268_), .B1(KEYINPUT70), .B2(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n277_), .A2(KEYINPUT70), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n205_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n211_), .A2(KEYINPUT12), .A3(new_n209_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n233_), .B2(new_n265_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n233_), .A2(KEYINPUT71), .A3(new_n265_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n259_), .B2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n287_), .A2(new_n277_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n258_), .A2(KEYINPUT8), .A3(new_n272_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n267_), .B1(new_n290_), .B2(new_n271_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n291_), .B2(new_n276_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n204_), .A3(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G120gat), .B(G148gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(G176gat), .B(G204gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n280_), .A2(new_n293_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(new_n280_), .B2(new_n293_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n202_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT13), .A3(new_n300_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G141gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G169gat), .B(G197gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G29gat), .B(G36gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G43gat), .B(G50gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G1gat), .A2(G8gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT14), .ZN(new_n315_));
  INV_X1    g114(.A(G15gat), .ZN(new_n316_));
  INV_X1    g115(.A(G22gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G15gat), .A2(G22gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n315_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n320_), .A2(KEYINPUT77), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n323_), .A2(KEYINPUT78), .A3(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G1gat), .B(G8gat), .Z(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT78), .B1(new_n323_), .B2(new_n324_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n326_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n313_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G229gat), .A2(G233gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n327_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n313_), .B(KEYINPUT15), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n328_), .A3(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n331_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n313_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n328_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n332_), .B1(new_n331_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n310_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n331_), .A2(new_n340_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n332_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n331_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n309_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n347_), .A3(KEYINPUT80), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(KEYINPUT22), .B(G169gat), .Z(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT81), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT82), .ZN(new_n361_));
  INV_X1    g160(.A(G183gat), .ZN(new_n362_));
  INV_X1    g161(.A(G190gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT23), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n361_), .B(new_n364_), .Z(new_n365_));
  NOR2_X1   g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n358_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT25), .B(G183gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n364_), .A2(new_n360_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n371_), .B(new_n372_), .C1(new_n357_), .C2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n367_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT83), .B(G15gat), .Z(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n375_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G127gat), .B(G134gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G120gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT85), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n380_), .A2(new_n381_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(KEYINPUT84), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n383_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n379_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389_));
  INV_X1    g188(.A(G43gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT30), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT31), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n388_), .B(new_n393_), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n397_), .B1(new_n402_), .B2(KEYINPUT1), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT87), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n400_), .A2(new_n401_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n403_), .A2(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n397_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n406_), .B2(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT87), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n412_), .B(KEYINPUT2), .ZN(new_n417_));
  NAND2_X1  g216(.A1(KEYINPUT88), .A2(KEYINPUT3), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(KEYINPUT88), .A2(KEYINPUT3), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n419_), .A2(new_n420_), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n414_), .A2(new_n418_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT89), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n421_), .A2(new_n417_), .A3(new_n425_), .A4(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n406_), .A2(new_n397_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT29), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT93), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G197gat), .B(G204gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G211gat), .B(G218gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT21), .ZN(new_n436_));
  OR4_X1    g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(G204gat), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n439_), .A2(G197gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT91), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n441_), .A3(KEYINPUT21), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(G197gat), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n440_), .B(new_n443_), .C1(KEYINPUT91), .C2(new_n436_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n444_), .A3(new_n435_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(KEYINPUT21), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n433_), .B1(new_n446_), .B2(new_n435_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n437_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT29), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(new_n416_), .B2(new_n429_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT93), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n432_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G228gat), .ZN(new_n454_));
  INV_X1    g253(.A(G233gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n431_), .A2(KEYINPUT90), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n448_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n458_), .B1(new_n431_), .B2(KEYINPUT90), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n453_), .A2(new_n456_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G78gat), .B(G106gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n396_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G50gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT28), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n430_), .B2(KEYINPUT29), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n411_), .A2(new_n415_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(KEYINPUT28), .A3(new_n449_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n466_), .A2(new_n317_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n317_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n464_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G22gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(new_n317_), .A3(new_n468_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(G50gat), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n457_), .A2(new_n459_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n431_), .A2(KEYINPUT93), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n456_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(new_n461_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n462_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n463_), .A2(new_n476_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n471_), .A2(new_n475_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n460_), .A2(new_n462_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n396_), .A4(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT4), .B1(new_n430_), .B2(new_n387_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n380_), .B(new_n381_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n416_), .A2(new_n429_), .A3(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n383_), .B(new_n385_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n467_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n494_), .B2(KEYINPUT4), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G225gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n430_), .A2(new_n387_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n499_), .B2(new_n492_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G1gat), .B(G29gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G85gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n502_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n500_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(new_n507_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G8gat), .B(G36gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT18), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G64gat), .B(G92gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n356_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n371_), .B1(new_n519_), .B2(new_n373_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n357_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(G176gat), .B2(new_n354_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n366_), .B1(new_n364_), .B2(new_n360_), .ZN(new_n523_));
  OAI22_X1  g322(.A1(new_n365_), .A2(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n448_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n525_), .B(KEYINPUT20), .C1(new_n375_), .C2(new_n448_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G226gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT19), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n375_), .A2(new_n448_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n524_), .A2(new_n448_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n529_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT20), .A4(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n527_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n518_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT96), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n526_), .A2(new_n529_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT95), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(new_n517_), .A3(new_n530_), .A4(new_n534_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT27), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT96), .B(new_n518_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT20), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n529_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(KEYINPUT98), .A3(new_n529_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT99), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n526_), .A2(new_n551_), .A3(new_n529_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n549_), .A2(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(KEYINPUT27), .B(new_n541_), .C1(new_n554_), .C2(new_n517_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n545_), .A2(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n489_), .A2(new_n513_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n517_), .A2(KEYINPUT32), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n540_), .A2(new_n558_), .A3(new_n530_), .A4(new_n534_), .ZN(new_n559_));
  OAI221_X1 g358(.A(new_n559_), .B1(new_n558_), .B2(new_n554_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n495_), .A2(new_n497_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n507_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n502_), .A2(new_n565_), .A3(new_n508_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT33), .B1(new_n510_), .B2(new_n507_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n560_), .A2(new_n569_), .B1(new_n488_), .B2(new_n484_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n395_), .B1(new_n557_), .B2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n545_), .A2(new_n555_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n489_), .A2(new_n572_), .A3(new_n512_), .A4(new_n394_), .ZN(new_n573_));
  AOI211_X1 g372(.A(new_n306_), .B(new_n353_), .C1(new_n571_), .C2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n580_));
  INV_X1    g379(.A(new_n285_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n283_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n275_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n580_), .B1(new_n583_), .B2(new_n336_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n291_), .B2(new_n313_), .ZN(new_n586_));
  AND4_X1   g385(.A1(new_n585_), .A2(new_n275_), .A3(new_n313_), .A4(new_n266_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n579_), .B(new_n584_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n275_), .A2(new_n313_), .A3(new_n266_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT74), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n275_), .A2(new_n585_), .A3(new_n313_), .A4(new_n266_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n579_), .B1(new_n593_), .B2(new_n584_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n578_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G190gat), .B(G218gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT36), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n584_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT73), .ZN(new_n601_));
  INV_X1    g400(.A(new_n578_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n588_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n595_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT75), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n595_), .B2(new_n603_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n575_), .B1(new_n604_), .B2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n589_), .A2(new_n594_), .A3(new_n578_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n602_), .B1(new_n601_), .B2(new_n588_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n607_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n599_), .B(KEYINPUT76), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n595_), .A2(new_n603_), .A3(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(KEYINPUT37), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n335_), .A2(new_n328_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n276_), .B(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT17), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n619_), .A2(new_n621_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n622_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n627_), .B(new_n628_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n622_), .B2(new_n630_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n617_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n574_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n574_), .A2(KEYINPUT100), .A3(new_n636_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(G1gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n513_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n643_), .A2(KEYINPUT101), .A3(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT101), .B1(new_n643_), .B2(new_n644_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n571_), .A2(new_n573_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n604_), .A2(new_n609_), .A3(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n595_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT103), .B1(new_n613_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n306_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n348_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n348_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT102), .B1(new_n306_), .B2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n634_), .A3(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n653_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n642_), .B1(new_n660_), .B2(new_n513_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n643_), .B1(new_n644_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n645_), .A2(new_n646_), .A3(new_n662_), .ZN(G1324gat));
  NOR2_X1   g462(.A1(new_n572_), .A2(G8gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n639_), .A2(new_n640_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n660_), .A2(new_n556_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G8gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT39), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n667_), .A2(KEYINPUT40), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  NAND3_X1  g474(.A1(new_n641_), .A2(new_n316_), .A3(new_n394_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT105), .Z(new_n677_));
  AOI21_X1  g476(.A(new_n316_), .B1(new_n660_), .B2(new_n394_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1326gat));
  AND2_X1   g479(.A1(new_n484_), .A2(new_n488_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n317_), .B1(new_n660_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n317_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT107), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n641_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n652_), .A2(new_n634_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n574_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n513_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n610_), .A2(new_n616_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(KEYINPUT108), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n560_), .A2(new_n569_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n489_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n572_), .A2(new_n512_), .A3(new_n488_), .A4(new_n484_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n394_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n573_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n617_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n696_), .A2(new_n704_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n656_), .A2(new_n635_), .A3(new_n658_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT108), .B(new_n693_), .C1(new_n647_), .C2(new_n617_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT43), .B1(new_n702_), .B2(new_n703_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT44), .B(new_n706_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT109), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n705_), .A2(new_n712_), .A3(KEYINPUT44), .A4(new_n706_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n707_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n513_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n692_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n714_), .B2(new_n556_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n556_), .B(KEYINPUT110), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT111), .B1(new_n690_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n574_), .A2(new_n724_), .A3(new_n689_), .A4(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n717_), .B1(new_n719_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n726_), .B(KEYINPUT45), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n705_), .A2(new_n706_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  AOI221_X4 g531(.A(new_n572_), .B1(new_n731_), .B2(new_n732_), .C1(new_n711_), .C2(new_n713_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n730_), .B(KEYINPUT46), .C1(new_n733_), .C2(new_n718_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n729_), .A2(new_n734_), .ZN(G1329gat));
  AOI21_X1  g534(.A(G43gat), .B1(new_n691_), .B2(new_n394_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n395_), .A2(new_n390_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n714_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n739_), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n736_), .B(new_n741_), .C1(new_n714_), .C2(new_n737_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1330gat));
  AOI21_X1  g542(.A(G50gat), .B1(new_n691_), .B2(new_n681_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n489_), .A2(new_n464_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n714_), .B2(new_n745_), .ZN(G1331gat));
  AND3_X1   g545(.A1(new_n350_), .A2(new_n634_), .A3(new_n351_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n653_), .A2(new_n654_), .A3(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(G57gat), .A3(new_n513_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT114), .ZN(new_n751_));
  INV_X1    g550(.A(G57gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n654_), .B(new_n348_), .C1(new_n571_), .C2(new_n573_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n636_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n512_), .B1(new_n754_), .B2(KEYINPUT113), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(KEYINPUT113), .B2(new_n754_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n751_), .B1(new_n752_), .B2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  INV_X1    g557(.A(new_n720_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n749_), .B2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT48), .Z(new_n761_));
  INV_X1    g560(.A(new_n754_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT115), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n761_), .A2(new_n766_), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n749_), .B2(new_n394_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT49), .Z(new_n771_));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n769_), .A3(new_n394_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1334gat));
  INV_X1    g572(.A(G78gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n749_), .B2(new_n681_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT50), .Z(new_n776_));
  NAND3_X1  g575(.A1(new_n762_), .A2(new_n774_), .A3(new_n681_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n753_), .A2(new_n689_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(G85gat), .A3(new_n512_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n306_), .A2(new_n657_), .A3(new_n635_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n705_), .A2(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n513_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n786_), .B2(new_n212_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT117), .ZN(G1336gat));
  OAI21_X1  g587(.A(new_n213_), .B1(new_n779_), .B2(new_n572_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT118), .Z(new_n790_));
  NOR2_X1   g589(.A1(new_n720_), .A2(new_n213_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n785_), .B2(new_n791_), .ZN(G1337gat));
  NOR3_X1   g591(.A1(new_n779_), .A2(new_n262_), .A3(new_n395_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n785_), .A2(new_n394_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n239_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g596(.A1(new_n779_), .A2(G106gat), .A3(new_n489_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n705_), .A2(new_n681_), .A3(new_n784_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G106gat), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT52), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n798_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n805_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n798_), .B(new_n807_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1339gat));
  NOR3_X1   g608(.A1(new_n681_), .A2(new_n556_), .A3(new_n395_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n304_), .A2(new_n300_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n338_), .A2(new_n341_), .A3(new_n310_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n309_), .B1(new_n343_), .B2(new_n332_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n331_), .A2(new_n344_), .A3(new_n337_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n811_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n300_), .A2(new_n348_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n276_), .B1(new_n275_), .B2(new_n266_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n287_), .B(new_n277_), .C1(new_n822_), .C2(KEYINPUT12), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n823_), .B2(new_n205_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n288_), .A2(KEYINPUT55), .A3(new_n204_), .A4(new_n292_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n205_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n298_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n298_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n820_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n819_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n820_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n831_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n298_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n833_), .B(new_n835_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n652_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n300_), .B(new_n818_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n843_), .A2(new_n842_), .B1(new_n610_), .B2(new_n616_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n840_), .A2(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n648_), .B1(new_n604_), .B2(new_n609_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n613_), .A2(KEYINPUT103), .A3(new_n650_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n850_), .A2(KEYINPUT121), .B1(new_n811_), .B2(new_n818_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n851_), .B2(new_n838_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT57), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n634_), .B1(new_n846_), .B2(new_n853_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n747_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n610_), .A3(new_n616_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT54), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n857_), .A3(new_n856_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n694_), .A2(KEYINPUT120), .A3(new_n855_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n857_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(KEYINPUT54), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n513_), .B(new_n810_), .C1(new_n854_), .C2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n348_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n845_), .A2(new_n844_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n852_), .B2(KEYINPUT57), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n840_), .A2(new_n841_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n635_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n858_), .B(new_n861_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n875_), .A2(KEYINPUT59), .A3(new_n513_), .A4(new_n810_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n353_), .B1(new_n869_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n867_), .B1(new_n877_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n865_), .B(new_n880_), .C1(KEYINPUT60), .C2(new_n879_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n654_), .B1(new_n869_), .B2(new_n876_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  OAI21_X1  g682(.A(G120gat), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  AOI211_X1 g683(.A(KEYINPUT123), .B(new_n654_), .C1(new_n869_), .C2(new_n876_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n881_), .B1(new_n884_), .B2(new_n885_), .ZN(G1341gat));
  INV_X1    g685(.A(G127gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n865_), .A2(new_n887_), .A3(new_n634_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n635_), .B1(new_n869_), .B2(new_n876_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n887_), .ZN(G1342gat));
  INV_X1    g689(.A(G134gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n865_), .A2(new_n891_), .A3(new_n849_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n694_), .B1(new_n869_), .B2(new_n876_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1343gat));
  AOI21_X1  g693(.A(new_n512_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n759_), .A2(new_n489_), .A3(new_n394_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n348_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n306_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n897_), .A2(new_n635_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  OAI21_X1  g704(.A(G162gat), .B1(new_n897_), .B2(new_n694_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n652_), .A2(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n897_), .B2(new_n907_), .ZN(G1347gat));
  NOR4_X1   g707(.A1(new_n720_), .A2(new_n513_), .A3(new_n681_), .A4(new_n395_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n875_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n348_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n911_), .A2(new_n912_), .A3(G169gat), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n911_), .A2(new_n354_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n911_), .B2(G169gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1348gat));
  NAND2_X1  g715(.A1(new_n910_), .A2(new_n306_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n634_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n369_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n362_), .B2(new_n919_), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n910_), .A2(new_n370_), .A3(new_n849_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n617_), .B(new_n909_), .C1(new_n854_), .C2(new_n863_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n923_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(KEYINPUT124), .B1(new_n923_), .B2(G190gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n922_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n922_), .B(new_n928_), .C1(new_n924_), .C2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1351gat));
  NAND3_X1  g729(.A1(new_n681_), .A2(new_n512_), .A3(new_n395_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n759_), .B1(new_n931_), .B2(KEYINPUT126), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n932_), .B1(KEYINPUT126), .B2(new_n931_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n875_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n657_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT127), .B(G197gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n934_), .A2(new_n654_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n439_), .ZN(G1353gat));
  INV_X1    g738(.A(new_n934_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n634_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  AND2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n941_), .B2(new_n942_), .ZN(G1354gat));
  OR3_X1    g744(.A1(new_n934_), .A2(G218gat), .A3(new_n652_), .ZN(new_n946_));
  OAI21_X1  g745(.A(G218gat), .B1(new_n934_), .B2(new_n694_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1355gat));
endmodule


