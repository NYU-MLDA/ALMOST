//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G134gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G232gat), .ZN(new_n207_));
  INV_X1    g006(.A(G233gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT67), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(KEYINPUT67), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(G99gat), .A4(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI211_X1 g025(.A(KEYINPUT8), .B(new_n212_), .C1(new_n222_), .C2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n213_), .A2(KEYINPUT68), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n216_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n213_), .A2(KEYINPUT68), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(G99gat), .A3(G106gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(KEYINPUT6), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n226_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n228_), .B1(new_n236_), .B2(new_n211_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n210_), .B1(new_n227_), .B2(new_n237_), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n215_), .A2(new_n217_), .A3(new_n213_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n219_), .A2(new_n220_), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n226_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n228_), .A3(new_n211_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n233_), .A2(new_n234_), .A3(KEYINPUT6), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT6), .B1(new_n233_), .B2(new_n234_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n212_), .B1(new_n245_), .B2(new_n226_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n242_), .B(KEYINPUT72), .C1(new_n246_), .C2(new_n228_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n238_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT9), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(G92gat), .ZN(new_n251_));
  INV_X1    g050(.A(G92gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT66), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  AOI22_X1  g053(.A1(KEYINPUT9), .A2(new_n211_), .B1(new_n254_), .B2(G85gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT10), .B(G99gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT64), .B(G106gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT65), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n255_), .B(new_n222_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n248_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT77), .B(G29gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G36gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G43gat), .B(G50gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n265_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT15), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n236_), .A2(new_n211_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT8), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n258_), .B(new_n259_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n255_), .A2(new_n222_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n272_), .A2(new_n242_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT78), .A3(new_n268_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n262_), .B1(new_n227_), .B2(new_n237_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n265_), .B(new_n266_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n270_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n209_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n209_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n270_), .A2(KEYINPUT79), .A3(new_n285_), .A4(new_n281_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n282_), .A2(KEYINPUT35), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n284_), .A2(new_n286_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n287_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT35), .B1(new_n295_), .B2(new_n289_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n202_), .B(new_n206_), .C1(new_n293_), .C2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n295_), .B(new_n289_), .C1(KEYINPUT35), .C2(new_n282_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT35), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n206_), .A2(new_n202_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n206_), .A2(new_n202_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT37), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n297_), .A2(KEYINPUT37), .A3(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G57gat), .A2(G64gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G57gat), .A2(G64gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G57gat), .ZN(new_n314_));
  INV_X1    g113(.A(G64gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT69), .B1(new_n316_), .B2(new_n309_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT11), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G71gat), .B(G78gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n312_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n316_), .A2(KEYINPUT69), .A3(new_n309_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT11), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT11), .B(new_n319_), .C1(new_n313_), .C2(new_n317_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G231gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G15gat), .B(G22gat), .Z(new_n330_));
  NAND2_X1  g129(.A1(G1gat), .A2(G8gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(KEYINPUT14), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT80), .ZN(new_n333_));
  XOR2_X1   g132(.A(G1gat), .B(G8gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n329_), .B(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G127gat), .B(G155gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(G183gat), .B(G211gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT17), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n342_), .A2(KEYINPUT81), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n336_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(KEYINPUT17), .B2(new_n341_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n348_), .B2(new_n336_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n308_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n335_), .B(new_n279_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G229gat), .A3(G233gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n335_), .A2(new_n279_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G229gat), .A2(G233gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n269_), .A2(new_n335_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G141gat), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G197gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n353_), .A2(new_n357_), .A3(new_n364_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT90), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT2), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n371_), .B(new_n373_), .C1(KEYINPUT90), .C2(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n370_), .ZN(new_n378_));
  OR3_X1    g177(.A1(new_n375_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(KEYINPUT1), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT89), .B1(new_n375_), .B2(KEYINPUT1), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n379_), .A2(new_n382_), .A3(new_n383_), .A4(new_n376_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n380_), .A2(new_n381_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n378_), .B(new_n372_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n377_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n388_), .A2(G113gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(G113gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G120gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(G120gat), .A3(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n387_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n377_), .A2(new_n394_), .A3(new_n393_), .A4(new_n386_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT99), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT99), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n387_), .A2(new_n400_), .A3(new_n395_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n396_), .A2(KEYINPUT4), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n401_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(KEYINPUT4), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n405_), .B2(new_n399_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G85gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(G1gat), .B(G29gat), .Z(new_n409_));
  XOR2_X1   g208(.A(new_n408_), .B(new_n409_), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n406_), .A2(new_n411_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G176gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n360_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT22), .B(G169gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n416_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT85), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(KEYINPUT85), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G183gat), .A2(G190gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT23), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n422_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(G183gat), .B2(G190gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n420_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT24), .B1(new_n360_), .B2(new_n416_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT25), .B(G183gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT26), .B(G190gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT24), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n422_), .A2(KEYINPUT23), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n424_), .B2(new_n422_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n432_), .A2(new_n435_), .A3(new_n437_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n427_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT86), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n427_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G211gat), .B(G218gat), .Z(new_n446_));
  XOR2_X1   g245(.A(G197gat), .B(G204gat), .Z(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT21), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT93), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT21), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n362_), .A2(G204gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n453_), .A2(new_n447_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n446_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n447_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n449_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n443_), .A2(new_n445_), .A3(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n460_), .A2(KEYINPUT20), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT19), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT96), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n432_), .A2(new_n425_), .A3(new_n435_), .A4(new_n437_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT97), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G183gat), .A2(G190gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n419_), .B1(new_n439_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT98), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n458_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(new_n464_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT103), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n445_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n444_), .B1(new_n427_), .B2(new_n441_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n458_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n465_), .A2(new_n468_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(KEYINPUT102), .Z(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT20), .B(new_n476_), .C1(new_n478_), .C2(new_n458_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n463_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n461_), .A2(KEYINPUT103), .A3(new_n464_), .A4(new_n470_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT18), .B(G64gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G92gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G8gat), .B(G36gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n461_), .A2(new_n470_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n464_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OR3_X1    g290(.A1(new_n466_), .A2(new_n458_), .A3(new_n469_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n463_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n492_), .A2(KEYINPUT20), .A3(new_n493_), .A4(new_n476_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n486_), .A3(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(KEYINPUT27), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497_));
  INV_X1    g296(.A(new_n495_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n486_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G78gat), .B(G106gat), .Z(new_n502_));
  OR3_X1    g301(.A1(new_n387_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT28), .B1(new_n387_), .B2(KEYINPUT29), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G22gat), .B(G50gat), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(G228gat), .A2(G233gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n377_), .B2(new_n386_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n459_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT94), .ZN(new_n516_));
  INV_X1    g315(.A(new_n514_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n512_), .B(KEYINPUT91), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n458_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n459_), .A2(new_n514_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(KEYINPUT94), .A3(new_n518_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(KEYINPUT95), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n515_), .A2(KEYINPUT94), .B1(new_n521_), .B2(new_n518_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n511_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n523_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n502_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n502_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n511_), .A2(new_n523_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n528_), .A2(new_n523_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(new_n533_), .C1(new_n534_), .C2(new_n511_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT30), .B(G43gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G227gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(G15gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G99gat), .Z(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n443_), .A2(new_n445_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n543_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n538_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n545_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n543_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n537_), .A3(new_n546_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(KEYINPUT87), .A3(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n395_), .B(KEYINPUT31), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n549_), .A2(new_n553_), .A3(KEYINPUT87), .A4(new_n555_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n536_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n558_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n501_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n412_), .A2(KEYINPUT33), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n406_), .A2(new_n565_), .A3(new_n411_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n404_), .A2(G225gat), .A3(G233gat), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n405_), .A2(KEYINPUT100), .A3(new_n399_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT100), .B1(new_n405_), .B2(new_n399_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n410_), .B(new_n568_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT101), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n405_), .A2(new_n399_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT100), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n405_), .A2(KEYINPUT100), .A3(new_n399_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n410_), .A4(new_n568_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n498_), .A2(new_n499_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n567_), .A2(new_n572_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n486_), .A2(KEYINPUT32), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n482_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n491_), .A2(new_n494_), .ZN(new_n584_));
  OAI221_X1 g383(.A(new_n583_), .B1(new_n584_), .B2(new_n582_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n561_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n536_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n415_), .A2(new_n563_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT75), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n325_), .A2(new_n326_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n272_), .A2(new_n242_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(new_n262_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT70), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n275_), .B2(new_n591_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n278_), .A2(KEYINPUT70), .A3(new_n327_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n594_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT71), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n591_), .B(new_n262_), .C1(new_n227_), .C2(new_n237_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT70), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n592_), .A2(new_n595_), .A3(new_n262_), .A4(new_n591_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n593_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT71), .B1(new_n606_), .B2(new_n600_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n600_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT73), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n603_), .A2(KEYINPUT73), .A3(new_n600_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n327_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n593_), .A2(KEYINPUT12), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT74), .B(G204gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT5), .B(G176gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n608_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n608_), .B2(new_n616_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT13), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n599_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n606_), .A2(KEYINPUT71), .A3(new_n600_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n616_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n621_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n608_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT13), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n590_), .B1(new_n626_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n625_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n630_), .A2(KEYINPUT13), .A3(new_n631_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(KEYINPUT75), .A3(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n351_), .A2(new_n367_), .A3(new_n589_), .A4(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G1gat), .A3(new_n415_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(new_n640_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n633_), .A2(new_n367_), .A3(new_n636_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT105), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n633_), .A2(new_n647_), .A3(new_n367_), .A4(new_n636_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(KEYINPUT106), .A3(new_n349_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n589_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n350_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n304_), .B1(new_n652_), .B2(KEYINPUT106), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n415_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n643_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n644_), .A2(new_n656_), .A3(new_n657_), .ZN(G1324gat));
  INV_X1    g457(.A(new_n501_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n651_), .A2(new_n653_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(G8gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT107), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n653_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n588_), .B1(new_n652_), .B2(KEYINPUT106), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n501_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(G8gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(KEYINPUT39), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n638_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n661_), .A3(new_n501_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT107), .B(new_n671_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n668_), .A2(KEYINPUT40), .A3(new_n670_), .A4(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  NAND3_X1  g476(.A1(new_n669_), .A2(new_n540_), .A3(new_n561_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n654_), .A2(new_n561_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n679_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT41), .B1(new_n679_), .B2(G15gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT108), .B(new_n678_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1326gat));
  INV_X1    g485(.A(G22gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n654_), .B2(new_n536_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT42), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n669_), .A2(new_n687_), .A3(new_n536_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(G29gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n588_), .A2(new_n304_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n645_), .A2(new_n349_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n692_), .B1(new_n695_), .B2(new_n415_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n581_), .A2(new_n585_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n559_), .A3(new_n587_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n562_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n561_), .B1(new_n531_), .B2(new_n535_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n415_), .B(new_n659_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n306_), .A2(new_n307_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  INV_X1    g504(.A(new_n307_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT37), .B1(new_n297_), .B2(new_n303_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT109), .B(new_n705_), .C1(new_n708_), .C2(new_n588_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n704_), .A2(new_n649_), .A3(new_n709_), .A4(new_n350_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G29gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n415_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n696_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT110), .B(new_n696_), .C1(new_n713_), .C2(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1328gat));
  NAND2_X1  g519(.A1(new_n712_), .A2(new_n501_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n710_), .A2(new_n711_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G36gat), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n693_), .A2(new_n724_), .A3(new_n501_), .A4(new_n694_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT45), .Z(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(KEYINPUT46), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n710_), .A2(new_n711_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n659_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n724_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n732_), .B2(new_n726_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n728_), .A2(new_n733_), .ZN(G1329gat));
  INV_X1    g533(.A(G43gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n695_), .B2(new_n559_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n712_), .A2(G43gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n561_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT47), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n741_), .B(new_n736_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1330gat));
  INV_X1    g542(.A(G50gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n695_), .B2(new_n587_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n712_), .A2(G50gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n536_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT111), .B(new_n745_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n588_), .A2(new_n367_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n637_), .A2(new_n350_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n304_), .A3(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n755_), .A2(new_n314_), .A3(new_n415_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n637_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n351_), .A2(new_n757_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n758_), .A2(KEYINPUT112), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(KEYINPUT112), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n753_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n714_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n756_), .B1(new_n762_), .B2(new_n314_), .ZN(G1332gat));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n315_), .A3(new_n501_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n755_), .A2(new_n659_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G64gat), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT113), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n768_), .A3(G64gat), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n767_), .A2(KEYINPUT48), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n767_), .B2(new_n769_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n764_), .B1(new_n770_), .B2(new_n771_), .ZN(G1333gat));
  NOR2_X1   g571(.A1(new_n559_), .A2(G71gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT114), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n761_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G71gat), .B1(new_n755_), .B2(new_n559_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT49), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1334gat));
  INV_X1    g577(.A(G78gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n761_), .A2(new_n779_), .A3(new_n536_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G78gat), .B1(new_n755_), .B2(new_n587_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT50), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n637_), .A2(new_n367_), .A3(new_n349_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n693_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n714_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n704_), .A2(new_n709_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n784_), .B(KEYINPUT115), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n714_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n789_), .B2(G85gat), .ZN(G1336gat));
  NAND2_X1  g589(.A1(new_n249_), .A2(G92gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n659_), .B1(new_n253_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n788_), .A3(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n785_), .A2(new_n501_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(G92gat), .B2(new_n794_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT116), .Z(G1337gat));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n561_), .A3(new_n788_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G99gat), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n559_), .A2(new_n256_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n785_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g601(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n704_), .A2(new_n788_), .A3(new_n709_), .A4(new_n536_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(G106gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT52), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n807_), .A3(G106gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n587_), .A2(new_n257_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n785_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n803_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n804_), .A2(new_n807_), .A3(G106gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n807_), .B1(new_n804_), .B2(G106gat), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n803_), .B(new_n811_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n812_), .A2(new_n816_), .ZN(G1339gat));
  NOR2_X1   g616(.A1(new_n501_), .A2(new_n415_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n366_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n352_), .A2(new_n355_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n354_), .A2(new_n356_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n821_), .B(new_n363_), .C1(new_n355_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n616_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n614_), .A2(new_n615_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n596_), .A2(new_n597_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n601_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n616_), .A2(new_n826_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n621_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n621_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n825_), .B(new_n631_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT58), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n308_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n367_), .A2(new_n631_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n833_), .A2(new_n834_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n623_), .A2(new_n624_), .ZN(new_n840_));
  OAI22_X1  g639(.A1(new_n838_), .A2(new_n839_), .B1(new_n840_), .B2(new_n824_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n304_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(KEYINPUT57), .A3(new_n304_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n350_), .B1(new_n837_), .B2(new_n846_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n367_), .A2(new_n626_), .A3(new_n632_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n306_), .A2(new_n349_), .A3(new_n307_), .A4(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT54), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n562_), .B(new_n819_), .C1(new_n847_), .C2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n367_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n850_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n699_), .A3(new_n818_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n562_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT118), .B1(new_n847_), .B2(new_n850_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n818_), .B(new_n859_), .C1(new_n860_), .C2(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n367_), .A2(G113gat), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT119), .Z(new_n864_));
  AOI21_X1  g663(.A(new_n852_), .B1(new_n862_), .B2(new_n864_), .ZN(G1340gat));
  OR2_X1    g664(.A1(new_n392_), .A2(KEYINPUT60), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n392_), .B1(new_n637_), .B2(KEYINPUT60), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n859_), .A2(new_n818_), .A3(new_n866_), .A4(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n851_), .A2(KEYINPUT120), .A3(new_n866_), .A4(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n637_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n392_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n851_), .B2(new_n349_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n350_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g676(.A(new_n304_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G134gat), .B1(new_n851_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n308_), .A2(G134gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT121), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n862_), .B2(new_n881_), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n853_), .A2(new_n700_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n367_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n883_), .A2(new_n884_), .A3(new_n819_), .ZN(new_n885_));
  INV_X1    g684(.A(G141gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1344gat));
  NOR3_X1   g686(.A1(new_n883_), .A2(new_n637_), .A3(new_n819_), .ZN(new_n888_));
  INV_X1    g687(.A(G148gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1345gat));
  AOI21_X1  g689(.A(new_n560_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n349_), .A3(new_n818_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT122), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n892_), .B(new_n894_), .ZN(G1346gat));
  NOR2_X1   g694(.A1(new_n883_), .A2(new_n819_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G162gat), .B1(new_n896_), .B2(new_n878_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n708_), .A2(new_n205_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n896_), .B2(new_n898_), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n659_), .A2(new_n714_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n367_), .A3(new_n561_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n418_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n853_), .A2(new_n587_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(KEYINPUT123), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n901_), .A2(KEYINPUT123), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n853_), .A2(new_n587_), .A3(new_n905_), .A4(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n907_), .A2(new_n908_), .A3(G169gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n907_), .B2(G169gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n904_), .B1(new_n909_), .B2(new_n910_), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n859_), .A2(new_n757_), .A3(new_n900_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G176gat), .ZN(G1349gat));
  AND2_X1   g712(.A1(new_n859_), .A2(new_n900_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n349_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(G183gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n349_), .A3(new_n433_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1350gat));
  NAND2_X1  g717(.A1(new_n914_), .A2(new_n308_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G190gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n878_), .A2(new_n434_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT124), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n914_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n923_), .ZN(G1351gat));
  NAND3_X1  g723(.A1(new_n891_), .A2(new_n367_), .A3(new_n900_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g725(.A1(new_n891_), .A2(new_n757_), .A3(new_n900_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n891_), .A2(new_n349_), .A3(new_n900_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT125), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT126), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n935_), .A2(KEYINPUT126), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n932_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT126), .B(new_n935_), .C1(new_n929_), .C2(new_n931_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1354gat));
  NAND3_X1  g739(.A1(new_n891_), .A2(new_n878_), .A3(new_n900_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT127), .ZN(new_n942_));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n891_), .A2(new_n944_), .A3(new_n878_), .A4(new_n900_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n943_), .A3(new_n945_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n891_), .A2(G218gat), .A3(new_n308_), .A4(new_n900_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1355gat));
endmodule


