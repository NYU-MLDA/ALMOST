//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_, new_n982_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211_));
  INV_X1    g010(.A(G155gat), .ZN(new_n212_));
  INV_X1    g011(.A(G162gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT84), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n210_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n214_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n209_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT86), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT86), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n229_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT85), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n225_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n205_), .B1(new_n224_), .B2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n208_), .A2(new_n209_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n222_), .A2(KEYINPUT84), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n219_), .A2(new_n220_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n231_), .A2(new_n233_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n227_), .A2(new_n228_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n235_), .A2(new_n236_), .ZN(new_n246_));
  NOR4_X1   g045(.A1(KEYINPUT85), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n244_), .B(new_n245_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n225_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n250_), .A3(new_n204_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n239_), .A2(KEYINPUT4), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n250_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n205_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G225gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G57gat), .B(G85gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT100), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(G1gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n263_));
  INV_X1    g062(.A(G29gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n262_), .B(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n258_), .B1(new_n239_), .B2(new_n251_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n262_), .A2(new_n265_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n262_), .A2(new_n265_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n257_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n267_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(KEYINPUT103), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT103), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n272_), .B(new_n276_), .C1(new_n273_), .C2(new_n267_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(KEYINPUT104), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT104), .B1(new_n275_), .B2(new_n277_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT80), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(G169gat), .A3(G176gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n290_), .B(new_n291_), .C1(G183gat), .C2(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(G169gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT22), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT24), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT81), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n290_), .A2(new_n291_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G190gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT26), .B1(new_n308_), .B2(KEYINPUT78), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT26), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(G183gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT25), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G183gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .A4(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n302_), .A2(KEYINPUT24), .A3(new_n303_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(new_n286_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n307_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n305_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n300_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G71gat), .B(G99gat), .ZN(new_n323_));
  INV_X1    g122(.A(G43gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n322_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(new_n205_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(G15gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT30), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT31), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n327_), .B(new_n332_), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n281_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n243_), .B2(new_n250_), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G197gat), .ZN(new_n338_));
  INV_X1    g137(.A(G197gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G204gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT21), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT90), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n338_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT21), .B1(new_n338_), .B2(new_n345_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT91), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n339_), .A2(G204gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n343_), .B1(new_n349_), .B2(KEYINPUT90), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT91), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n338_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n342_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n343_), .B2(new_n341_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n344_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n358_), .A2(KEYINPUT92), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(KEYINPUT92), .ZN(new_n360_));
  OAI22_X1  g159(.A1(new_n336_), .A2(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT91), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n351_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n356_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n344_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n360_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n223_), .A2(new_n220_), .A3(new_n219_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n368_), .A2(new_n240_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n366_), .B(new_n367_), .C1(new_n335_), .C2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT95), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT95), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n361_), .A2(new_n370_), .A3(new_n375_), .A4(new_n372_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G22gat), .B(G50gat), .Z(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n369_), .B2(new_n335_), .ZN(new_n380_));
  AND4_X1   g179(.A1(new_n335_), .A2(new_n243_), .A3(new_n250_), .A4(new_n379_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n377_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(new_n253_), .B2(KEYINPUT29), .ZN(new_n384_));
  INV_X1    g183(.A(new_n377_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n369_), .A2(new_n335_), .A3(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n382_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n383_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n374_), .B(new_n376_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n361_), .A2(new_n370_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n372_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n361_), .A2(new_n370_), .A3(KEYINPUT93), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(KEYINPUT94), .A3(new_n394_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n390_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n389_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n391_), .A2(new_n371_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n373_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n382_), .A2(new_n387_), .A3(new_n383_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n408_), .B(new_n409_), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n322_), .B2(new_n357_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT97), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n294_), .A2(new_n296_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n286_), .B1(new_n417_), .B2(new_n297_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT98), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n292_), .B(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422_));
  INV_X1    g221(.A(new_n303_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n306_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT96), .B1(new_n304_), .B2(new_n306_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n318_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n314_), .A2(new_n316_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT26), .B(G190gat), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n431_), .A2(new_n282_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n421_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n366_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT19), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n413_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n418_), .A2(new_n420_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n412_), .B1(new_n442_), .B2(new_n357_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n319_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT81), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n321_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n299_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n366_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n440_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT102), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n441_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  AOI211_X1 g250(.A(KEYINPUT102), .B(new_n440_), .C1(new_n443_), .C2(new_n448_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n411_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT20), .B1(new_n447_), .B2(new_n366_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n442_), .A2(new_n357_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n439_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n443_), .A2(new_n440_), .A3(new_n448_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n410_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(KEYINPUT27), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n357_), .A2(new_n421_), .A3(new_n435_), .ZN(new_n460_));
  AND4_X1   g259(.A1(KEYINPUT20), .A2(new_n448_), .A3(new_n440_), .A4(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n440_), .B1(new_n413_), .B2(new_n437_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n411_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n458_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT27), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n453_), .A2(new_n459_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n406_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n334_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n399_), .B2(new_n405_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n275_), .A2(new_n277_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT104), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n278_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT105), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n333_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n410_), .A2(KEYINPUT32), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n456_), .A2(new_n457_), .A3(new_n477_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n275_), .A3(new_n277_), .A4(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n272_), .B(KEYINPUT33), .C1(new_n273_), .C2(new_n267_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT101), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n274_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n239_), .A2(new_n258_), .A3(new_n251_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n266_), .B(new_n486_), .C1(new_n258_), .C2(new_n256_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n485_), .A2(new_n458_), .A3(new_n463_), .A4(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n406_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n391_), .A2(new_n392_), .ZN(new_n491_));
  AND4_X1   g290(.A1(KEYINPUT94), .A2(new_n491_), .A3(new_n371_), .A4(new_n394_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT94), .B1(new_n393_), .B2(new_n394_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n404_), .B1(new_n494_), .B2(new_n390_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n495_), .A2(new_n278_), .A3(new_n472_), .A4(new_n466_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n490_), .A2(new_n496_), .A3(KEYINPUT105), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n468_), .B1(new_n476_), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT69), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n499_), .A2(KEYINPUT69), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(KEYINPUT69), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508_));
  INV_X1    g307(.A(G1gat), .ZN(new_n509_));
  INV_X1    g308(.A(G8gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT14), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G1gat), .B(G8gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n503_), .A2(new_n514_), .A3(new_n506_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT75), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n519_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n516_), .A2(new_n520_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n507_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n503_), .A2(new_n506_), .A3(new_n527_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n514_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT76), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n529_), .A2(new_n533_), .A3(new_n530_), .A4(new_n514_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n526_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT77), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n525_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n523_), .A2(new_n524_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n540_), .B1(new_n543_), .B2(new_n535_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT10), .B(G99gat), .Z(new_n549_));
  INV_X1    g348(.A(G106gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G85gat), .B(G92gat), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT9), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554_));
  INV_X1    g353(.A(G85gat), .ZN(new_n555_));
  INV_X1    g354(.A(G92gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT6), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(G99gat), .A3(G106gat), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n554_), .A2(new_n557_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n551_), .A2(new_n553_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT64), .ZN(new_n564_));
  NOR2_X1   g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT7), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n559_), .A2(new_n561_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n552_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT8), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G57gat), .B(G64gat), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n571_), .A2(KEYINPUT11), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(KEYINPUT11), .ZN(new_n573_));
  XOR2_X1   g372(.A(G71gat), .B(G78gat), .Z(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n564_), .A2(new_n570_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT65), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT64), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n563_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT8), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n569_), .B(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n577_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n548_), .B1(new_n580_), .B2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n548_), .B1(new_n585_), .B2(new_n577_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n585_), .A2(KEYINPUT12), .A3(new_n577_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n564_), .A2(new_n570_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n577_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n588_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT66), .B(KEYINPUT5), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT67), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n595_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n587_), .A2(new_n594_), .A3(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT13), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(KEYINPUT13), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n564_), .A2(new_n570_), .A3(new_n507_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT35), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT71), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(KEYINPUT35), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n529_), .A2(new_n530_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n611_), .B(new_n618_), .C1(new_n585_), .C2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT71), .A3(new_n615_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n591_), .A2(new_n530_), .A3(new_n529_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n615_), .A2(KEYINPUT71), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n611_), .A4(new_n618_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT36), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n621_), .A2(new_n624_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n627_), .A2(KEYINPUT36), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT72), .B(new_n634_), .C1(new_n621_), .C2(new_n624_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n629_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT37), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n514_), .B(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(new_n592_), .ZN(new_n640_));
  XOR2_X1   g439(.A(G127gat), .B(G155gat), .Z(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT16), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT17), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT73), .Z(new_n648_));
  AND2_X1   g447(.A1(new_n644_), .A2(new_n645_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n640_), .A2(new_n646_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT74), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n610_), .A2(new_n637_), .A3(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n498_), .A2(new_n546_), .A3(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n509_), .A3(new_n473_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT38), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n609_), .A2(new_n546_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n651_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n334_), .A2(new_n467_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n490_), .A2(new_n496_), .A3(KEYINPUT105), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n281_), .A2(new_n475_), .A3(new_n495_), .A4(new_n466_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n333_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n662_), .B1(new_n668_), .B2(new_n636_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n636_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT105), .B1(new_n469_), .B2(new_n473_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n482_), .B(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n464_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n485_), .A4(new_n487_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n495_), .B1(new_n675_), .B2(new_n481_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n666_), .B(new_n665_), .C1(new_n671_), .C2(new_n676_), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT106), .B(new_n670_), .C1(new_n677_), .C2(new_n663_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n661_), .B1(new_n669_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT106), .B1(new_n498_), .B2(new_n670_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n668_), .A2(new_n662_), .A3(new_n636_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(KEYINPUT107), .A3(new_n661_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n281_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n657_), .B1(new_n686_), .B2(new_n509_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT108), .Z(G1324gat));
  OAI21_X1  g487(.A(G8gat), .B1(new_n679_), .B2(new_n466_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n689_), .A2(KEYINPUT39), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(KEYINPUT39), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n466_), .A2(G8gat), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n690_), .A2(new_n691_), .B1(new_n655_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n693_), .B(new_n695_), .ZN(G1325gat));
  AOI21_X1  g495(.A(new_n666_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT110), .B1(new_n697_), .B2(new_n329_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT107), .B1(new_n684_), .B2(new_n661_), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n680_), .B(new_n660_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n333_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(G15gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n698_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n655_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n698_), .A2(KEYINPUT41), .A3(new_n703_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(G1326gat));
  INV_X1    g508(.A(G22gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n655_), .A2(new_n710_), .A3(new_n495_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n406_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n712_), .A2(KEYINPUT42), .A3(new_n710_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n495_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G22gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n713_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT111), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n719_), .B(new_n711_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1327gat));
  NOR2_X1   g520(.A1(new_n498_), .A2(new_n546_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n651_), .B(KEYINPUT74), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n670_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n609_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n264_), .A3(new_n473_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n498_), .A2(new_n637_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT37), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n636_), .B(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n668_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT43), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n658_), .A2(new_n723_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n730_), .B2(new_n734_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT112), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n281_), .B1(new_n741_), .B2(KEYINPUT44), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G29gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n744_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n727_), .B1(new_n747_), .B2(new_n748_), .ZN(G1328gat));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750_));
  INV_X1    g549(.A(G36gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n741_), .A2(KEYINPUT44), .ZN(new_n752_));
  INV_X1    g551(.A(new_n466_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n743_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n466_), .B(KEYINPUT114), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n726_), .A2(new_n751_), .A3(new_n758_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT45), .Z(new_n760_));
  OAI21_X1  g559(.A(new_n750_), .B1(new_n756_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n760_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n754_), .B1(new_n742_), .B2(new_n740_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n762_), .B(KEYINPUT46), .C1(new_n751_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1329gat));
  NOR2_X1   g564(.A1(new_n666_), .A2(new_n324_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n742_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n741_), .B2(KEYINPUT112), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n752_), .B(new_n766_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n726_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n324_), .B1(new_n771_), .B2(new_n666_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(G1330gat));
  AOI21_X1  g574(.A(G50gat), .B1(new_n726_), .B2(new_n495_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n743_), .A2(new_n752_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n495_), .A2(G50gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(G1331gat));
  NOR2_X1   g578(.A1(new_n610_), .A2(new_n545_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n684_), .A2(new_n653_), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G57gat), .B1(new_n781_), .B2(new_n281_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n732_), .A2(new_n723_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n609_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT116), .Z(new_n785_));
  NOR2_X1   g584(.A1(new_n498_), .A2(new_n545_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n281_), .A2(G57gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n782_), .B1(new_n787_), .B2(new_n788_), .ZN(G1332gat));
  OR3_X1    g588(.A1(new_n787_), .A2(G64gat), .A3(new_n757_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G64gat), .B1(new_n781_), .B2(new_n757_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT48), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(KEYINPUT48), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(G1333gat));
  OR3_X1    g593(.A1(new_n787_), .A2(G71gat), .A3(new_n666_), .ZN(new_n795_));
  OAI21_X1  g594(.A(G71gat), .B1(new_n781_), .B2(new_n666_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(KEYINPUT49), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(KEYINPUT49), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n795_), .B1(new_n797_), .B2(new_n798_), .ZN(G1334gat));
  OR3_X1    g598(.A1(new_n787_), .A2(G78gat), .A3(new_n406_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G78gat), .B1(new_n781_), .B2(new_n406_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(KEYINPUT50), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(KEYINPUT50), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n800_), .B1(new_n802_), .B2(new_n803_), .ZN(G1335gat));
  NOR2_X1   g603(.A1(new_n724_), .A2(new_n610_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n786_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n555_), .A3(new_n473_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n735_), .A2(new_n723_), .A3(new_n780_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n473_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n810_), .B2(new_n555_), .ZN(G1336gat));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n556_), .A3(new_n753_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n809_), .A2(new_n758_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n556_), .ZN(G1337gat));
  AND3_X1   g613(.A1(new_n807_), .A2(new_n333_), .A3(new_n549_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n809_), .A2(new_n333_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(G99gat), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g617(.A1(new_n807_), .A2(new_n550_), .A3(new_n495_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n735_), .A2(new_n495_), .A3(new_n723_), .A4(new_n780_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(G106gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(G106gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g624(.A1(new_n589_), .A2(new_n593_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n548_), .B1(new_n826_), .B2(new_n580_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT55), .B(new_n588_), .C1(new_n589_), .C2(new_n593_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n594_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n602_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(KEYINPUT56), .A3(new_n602_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n539_), .B1(new_n543_), .B2(new_n535_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n516_), .A2(new_n521_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n840_), .B2(new_n539_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n604_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT58), .B1(new_n836_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT118), .B1(new_n844_), .B2(new_n637_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT58), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n732_), .B(new_n848_), .C1(new_n846_), .C2(KEYINPUT58), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n845_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n545_), .A2(KEYINPUT117), .A3(new_n604_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT117), .B1(new_n545_), .B2(new_n604_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n855_), .A2(new_n836_), .B1(new_n605_), .B2(new_n841_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n856_), .B2(new_n670_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n541_), .B1(new_n525_), .B2(new_n536_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n543_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n604_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n831_), .A2(KEYINPUT56), .A3(new_n602_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n602_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n862_), .B(new_n852_), .C1(new_n863_), .C2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n605_), .A2(new_n841_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT57), .A3(new_n636_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n857_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n723_), .B1(new_n850_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT54), .B1(new_n654_), .B2(new_n545_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n783_), .A2(new_n874_), .A3(new_n546_), .A4(new_n610_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n867_), .B2(new_n636_), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n851_), .B(new_n670_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n845_), .A2(new_n849_), .A3(new_n847_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n653_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT119), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n872_), .A2(new_n876_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n473_), .A2(new_n333_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n467_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(KEYINPUT59), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n659_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n873_), .A2(new_n875_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n883_), .A2(new_n887_), .B1(KEYINPUT59), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G113gat), .B1(new_n892_), .B2(new_n546_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n546_), .A2(G113gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n890_), .B2(new_n894_), .ZN(G1340gat));
  XNOR2_X1  g694(.A(KEYINPUT120), .B(G120gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT60), .B1(new_n609_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n609_), .B1(new_n890_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n891_), .B2(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n890_), .A2(KEYINPUT60), .A3(new_n897_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT121), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  INV_X1    g702(.A(new_n901_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n887_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n889_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n882_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n890_), .A2(KEYINPUT59), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n898_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n903_), .B(new_n904_), .C1(new_n909_), .C2(new_n896_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n902_), .A2(new_n910_), .ZN(G1341gat));
  OAI21_X1  g710(.A(G127gat), .B1(new_n892_), .B2(new_n651_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n723_), .A2(G127gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n890_), .B2(new_n913_), .ZN(G1342gat));
  NOR2_X1   g713(.A1(new_n890_), .A2(new_n636_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(G134gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n732_), .A2(G134gat), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT122), .Z(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n891_), .B2(new_n918_), .ZN(G1343gat));
  OAI21_X1  g718(.A(new_n651_), .B1(new_n850_), .B2(new_n869_), .ZN(new_n920_));
  AOI211_X1 g719(.A(new_n406_), .B(new_n333_), .C1(new_n920_), .C2(new_n876_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n473_), .A3(new_n757_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n546_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT123), .B(G141gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1344gat));
  NOR2_X1   g724(.A1(new_n922_), .A2(new_n610_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT124), .B(G148gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1345gat));
  NOR2_X1   g727(.A1(new_n922_), .A2(new_n723_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT61), .B(G155gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n922_), .B2(new_n637_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n670_), .A2(new_n213_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n922_), .B2(new_n933_), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n757_), .A2(new_n334_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n495_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n876_), .B1(new_n881_), .B2(KEYINPUT119), .ZN(new_n938_));
  AOI211_X1 g737(.A(new_n871_), .B(new_n653_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940_), .B2(new_n546_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n941_), .A2(KEYINPUT62), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(KEYINPUT62), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n883_), .A2(KEYINPUT125), .A3(new_n937_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n545_), .A2(new_n417_), .ZN(new_n950_));
  OAI22_X1  g749(.A1(new_n942_), .A2(new_n943_), .B1(new_n949_), .B2(new_n950_), .ZN(G1348gat));
  OAI21_X1  g750(.A(new_n609_), .B1(new_n946_), .B2(new_n948_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n495_), .B1(new_n920_), .B2(new_n876_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n936_), .A2(new_n297_), .A3(new_n610_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n952_), .A2(new_n297_), .B1(new_n953_), .B2(new_n954_), .ZN(G1349gat));
  NAND3_X1  g754(.A1(new_n953_), .A2(new_n653_), .A3(new_n935_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n313_), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n651_), .A2(new_n432_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n959_), .B2(KEYINPUT126), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961_));
  AOI211_X1 g760(.A(new_n961_), .B(new_n958_), .C1(new_n945_), .C2(new_n947_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n960_), .A2(new_n962_), .ZN(G1350gat));
  NAND2_X1  g762(.A1(new_n670_), .A2(new_n433_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n637_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n965_));
  OAI22_X1  g764(.A1(new_n949_), .A2(new_n964_), .B1(new_n965_), .B2(new_n308_), .ZN(G1351gat));
  NOR2_X1   g765(.A1(new_n757_), .A2(new_n473_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n921_), .A2(new_n967_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n968_), .A2(new_n546_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(new_n339_), .ZN(G1352gat));
  NOR2_X1   g769(.A1(new_n968_), .A2(new_n610_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(new_n337_), .ZN(G1353gat));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  AND2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  NOR4_X1   g773(.A1(new_n968_), .A2(new_n651_), .A3(new_n973_), .A4(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n968_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(new_n659_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n975_), .B1(new_n977_), .B2(new_n973_), .ZN(G1354gat));
  AND3_X1   g777(.A1(new_n976_), .A2(G218gat), .A3(new_n732_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n968_), .A2(KEYINPUT127), .A3(new_n636_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n980_), .A2(G218gat), .ZN(new_n981_));
  OAI21_X1  g780(.A(KEYINPUT127), .B1(new_n968_), .B2(new_n636_), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n979_), .B1(new_n981_), .B2(new_n982_), .ZN(G1355gat));
endmodule


