//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT2), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT87), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .A4(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(new_n209_), .B2(KEYINPUT87), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n203_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216_));
  OR3_X1    g015(.A1(new_n212_), .A2(new_n216_), .A3(KEYINPUT1), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n214_), .B1(KEYINPUT1), .B2(new_n212_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G141gat), .B(G148gat), .Z(new_n221_));
  AOI22_X1  g020(.A1(new_n211_), .A2(new_n215_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G22gat), .B(G50gat), .Z(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT95), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G204gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G197gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT21), .B1(new_n237_), .B2(KEYINPUT90), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G204gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n241_), .B2(KEYINPUT90), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n240_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(KEYINPUT21), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n247_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n248_), .A2(KEYINPUT21), .A3(new_n244_), .A4(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT92), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n246_), .A2(KEYINPUT92), .A3(new_n250_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G233gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n256_), .A2(KEYINPUT89), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(KEYINPUT89), .ZN(new_n258_));
  OAI21_X1  g057(.A(G228gat), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(KEYINPUT93), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT93), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n254_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n259_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n251_), .A2(KEYINPUT94), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT94), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n246_), .A2(new_n269_), .A3(new_n250_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n222_), .A2(new_n223_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n267_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G78gat), .B(G106gat), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n266_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n266_), .B2(new_n273_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n235_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n265_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n264_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n273_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n274_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n266_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n234_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT18), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT23), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G190gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT25), .B(G183gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(KEYINPUT24), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n307_), .A2(KEYINPUT97), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(KEYINPUT97), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n296_), .B(new_n300_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n299_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n305_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(KEYINPUT98), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(KEYINPUT98), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n295_), .A2(KEYINPUT80), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n295_), .A2(KEYINPUT80), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n293_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n314_), .A2(new_n315_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n268_), .A2(new_n310_), .A3(new_n320_), .A4(new_n270_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n305_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT78), .B(G183gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n292_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n296_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G169gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(G176gat), .B1(new_n327_), .B2(KEYINPUT82), .ZN(new_n328_));
  XOR2_X1   g127(.A(KEYINPUT81), .B(G169gat), .Z(new_n329_));
  OAI221_X1 g128(.A(new_n328_), .B1(KEYINPUT82), .B2(new_n327_), .C1(new_n329_), .C2(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n295_), .B(KEYINPUT80), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n294_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n291_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n323_), .B2(new_n334_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n322_), .A2(new_n297_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n336_), .A2(new_n301_), .B1(new_n304_), .B2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n333_), .B(new_n300_), .C1(new_n338_), .C2(KEYINPUT79), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(KEYINPUT79), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n331_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n321_), .B(KEYINPUT20), .C1(new_n342_), .C2(new_n264_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n264_), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n345_), .B(KEYINPUT96), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n310_), .A2(new_n320_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n351_), .B2(new_n251_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n290_), .B1(new_n346_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n255_), .B2(new_n341_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT99), .B1(new_n351_), .B2(new_n251_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n251_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT99), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n357_), .A2(new_n310_), .A3(new_n358_), .A4(new_n320_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n345_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n347_), .A2(new_n352_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n348_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n354_), .B1(new_n365_), .B2(new_n290_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G85gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G57gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT85), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(KEYINPUT85), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n373_), .B(KEYINPUT85), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI211_X1 g179(.A(KEYINPUT4), .B(new_n222_), .C1(new_n377_), .C2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n377_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n211_), .A2(new_n215_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n220_), .A2(new_n221_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT100), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n222_), .A2(new_n380_), .A3(KEYINPUT100), .A4(new_n377_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI211_X1 g188(.A(new_n372_), .B(new_n381_), .C1(new_n389_), .C2(KEYINPUT4), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n372_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n371_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n381_), .B1(new_n389_), .B2(KEYINPUT4), .ZN(new_n394_));
  INV_X1    g193(.A(new_n372_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n370_), .A3(new_n391_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n366_), .A2(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n362_), .A2(new_n364_), .A3(new_n289_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n289_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n394_), .A2(new_n372_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n370_), .B1(new_n389_), .B2(new_n395_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n402_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n397_), .A2(new_n403_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n285_), .B(new_n399_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n393_), .A2(new_n397_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n346_), .A2(new_n353_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n289_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n362_), .A2(new_n364_), .A3(new_n289_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT27), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n411_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n285_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G43gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(G15gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n423_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n341_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n382_), .B(KEYINPUT31), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n431_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n429_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n341_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT84), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n433_), .B(new_n434_), .C1(new_n439_), .C2(new_n427_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n434_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n427_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n442_), .B2(new_n432_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n410_), .A2(new_n421_), .A3(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n285_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n444_), .A2(new_n398_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT101), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n285_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n411_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT101), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n445_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G43gat), .B(G50gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT69), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n456_), .A2(KEYINPUT69), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n455_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n456_), .A2(KEYINPUT69), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n457_), .A3(new_n454_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n460_), .A2(KEYINPUT15), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT15), .B1(new_n460_), .B2(new_n462_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT74), .B(G8gat), .ZN(new_n466_));
  INV_X1    g265(.A(G1gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G8gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n465_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT76), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n460_), .A2(new_n462_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n475_), .B(new_n481_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n478_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n477_), .A2(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT77), .ZN(new_n487_));
  XOR2_X1   g286(.A(G169gat), .B(G197gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n485_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n494_));
  XOR2_X1   g293(.A(G71gat), .B(G78gat), .Z(new_n495_));
  OR2_X1    g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n495_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT8), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  INV_X1    g307(.A(G99gat), .ZN(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n502_), .B1(new_n507_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT65), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(new_n502_), .C1(new_n507_), .C2(new_n513_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n500_), .A2(new_n501_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(new_n513_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n504_), .A2(new_n506_), .A3(new_n520_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n519_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n515_), .B(new_n517_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT10), .B(G99gat), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n510_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT64), .B(G92gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(G85gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n518_), .A2(KEYINPUT9), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n504_), .A2(new_n506_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n499_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n492_), .B1(new_n535_), .B2(KEYINPUT12), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n515_), .A2(new_n517_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n511_), .A2(new_n512_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n523_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n525_), .B1(new_n540_), .B2(new_n518_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n534_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n499_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT68), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n536_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(KEYINPUT12), .A3(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT67), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT67), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n542_), .A2(new_n550_), .A3(KEYINPUT12), .A4(new_n543_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n542_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n499_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n547_), .A2(new_n552_), .A3(new_n553_), .A4(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n553_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n555_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n535_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n556_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n491_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n556_), .A2(new_n559_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n556_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(KEYINPUT13), .A3(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n499_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n475_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(KEYINPUT17), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n578_), .B1(new_n582_), .B2(new_n576_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  INV_X1    g386(.A(new_n481_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT70), .B1(new_n542_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n526_), .A2(new_n590_), .A3(new_n481_), .A4(new_n534_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT34), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n465_), .A2(new_n542_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n592_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n596_), .A2(new_n593_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(KEYINPUT71), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n592_), .A2(new_n603_), .A3(new_n599_), .A4(new_n597_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT72), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT36), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n587_), .B1(new_n613_), .B2(KEYINPUT73), .ZN(new_n614_));
  INV_X1    g413(.A(new_n611_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n616_));
  AOI211_X1 g415(.A(new_n601_), .B(new_n604_), .C1(new_n592_), .C2(new_n597_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n607_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n613_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n619_), .B(new_n613_), .C1(KEYINPUT73), .C2(new_n587_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n586_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n453_), .A2(new_n490_), .A3(new_n572_), .A4(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT102), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n411_), .A2(G1gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT103), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT103), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n446_), .A2(KEYINPUT101), .A3(new_n447_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n451_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n440_), .A2(new_n443_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n634_), .A2(new_n635_), .B1(new_n637_), .B2(new_n410_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n620_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n572_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n490_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n586_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n411_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n633_), .A2(new_n648_), .A3(new_n649_), .ZN(G1324gat));
  NAND2_X1  g449(.A1(new_n413_), .A2(new_n418_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G8gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT39), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n625_), .A2(new_n651_), .A3(new_n466_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n636_), .A2(new_n425_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n624_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n425_), .B1(new_n646_), .B2(new_n636_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  OAI21_X1  g465(.A(G22gat), .B1(new_n647_), .B2(new_n285_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT42), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n285_), .A2(G22gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n624_), .B2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n620_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n572_), .A2(new_n586_), .A3(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n638_), .A2(new_n644_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G29gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n398_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  INV_X1    g476(.A(new_n586_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n643_), .A2(new_n678_), .A3(new_n644_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n621_), .A2(new_n622_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT108), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n638_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n453_), .A2(new_n684_), .A3(new_n681_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n680_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n677_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n621_), .A2(new_n622_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT108), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n684_), .B1(new_n453_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n681_), .A2(new_n684_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n638_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n679_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(KEYINPUT109), .A3(new_n694_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n687_), .A2(new_n695_), .B1(KEYINPUT44), .B2(new_n686_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n398_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n676_), .B1(new_n697_), .B2(G29gat), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT110), .B(new_n674_), .C1(new_n696_), .C2(new_n398_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n675_), .B1(new_n698_), .B2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n687_), .A2(new_n695_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n686_), .A2(KEYINPUT44), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n651_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(G36gat), .B1(new_n413_), .B2(new_n418_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n673_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT45), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n673_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n711_), .A2(new_n713_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n704_), .B1(new_n708_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n714_), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n703_), .B(new_n716_), .C1(new_n707_), .C2(G36gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1329gat));
  NAND3_X1  g517(.A1(new_n696_), .A2(G43gat), .A3(new_n636_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT112), .B(G43gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n673_), .B2(new_n636_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n719_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n673_), .B2(new_n420_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n420_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n696_), .B2(new_n729_), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n638_), .A2(new_n490_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n731_), .A2(new_n643_), .A3(new_n623_), .ZN(new_n732_));
  INV_X1    g531(.A(G57gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n398_), .ZN(new_n734_));
  AND4_X1   g533(.A1(new_n644_), .A2(new_n642_), .A3(new_n643_), .A4(new_n678_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n398_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n736_), .B2(new_n733_), .ZN(G1332gat));
  INV_X1    g536(.A(G64gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n735_), .B2(new_n651_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n732_), .A2(new_n738_), .A3(new_n651_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n735_), .B2(new_n636_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT49), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n732_), .A2(new_n744_), .A3(new_n636_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1334gat));
  INV_X1    g547(.A(G78gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n735_), .B2(new_n420_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT50), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n732_), .A2(new_n749_), .A3(new_n420_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1335gat));
  NAND3_X1  g552(.A1(new_n643_), .A2(new_n644_), .A3(new_n586_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n411_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n572_), .A2(new_n678_), .A3(new_n620_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n731_), .A2(new_n758_), .ZN(new_n759_));
  OR3_X1    g558(.A1(new_n759_), .A2(G85gat), .A3(new_n411_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1336gat));
  INV_X1    g560(.A(new_n759_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G92gat), .B1(new_n762_), .B2(new_n651_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n651_), .A2(new_n529_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n755_), .B2(new_n764_), .ZN(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n756_), .B2(new_n444_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n636_), .A2(new_n527_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n759_), .B2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g568(.A1(new_n762_), .A2(new_n510_), .A3(new_n420_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n771_));
  INV_X1    g570(.A(new_n754_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n420_), .B(new_n772_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G106gat), .B1(new_n773_), .B2(KEYINPUT114), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n755_), .B2(new_n420_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n771_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n771_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n774_), .A2(new_n777_), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n770_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n770_), .B(new_n783_), .C1(new_n779_), .C2(new_n781_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1339gat));
  NOR3_X1   g586(.A1(new_n449_), .A2(new_n411_), .A3(new_n444_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n557_), .B2(KEYINPUT118), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n550_), .B1(new_n535_), .B2(KEYINPUT12), .ZN(new_n792_));
  INV_X1    g591(.A(new_n551_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n555_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT68), .B1(new_n544_), .B2(new_n545_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n492_), .B(KEYINPUT12), .C1(new_n542_), .C2(new_n543_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n791_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n791_), .B1(new_n790_), .B2(new_n557_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n547_), .A2(new_n552_), .A3(new_n555_), .A4(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n563_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n563_), .A4(new_n800_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n804_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n547_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n564_), .B1(new_n808_), .B2(new_n791_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n800_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n565_), .A2(new_n644_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n477_), .B(new_n480_), .C1(new_n476_), .C2(new_n588_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n489_), .B1(new_n483_), .B2(new_n479_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n485_), .A2(new_n489_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n671_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n570_), .A2(new_n816_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT121), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n570_), .A2(new_n821_), .A3(new_n816_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n805_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n820_), .B(new_n822_), .C1(new_n810_), .C2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n688_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n803_), .A2(new_n805_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n820_), .A4(new_n822_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n818_), .A2(KEYINPUT57), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n830_));
  OAI21_X1  g629(.A(new_n812_), .B1(new_n807_), .B2(new_n810_), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n804_), .B(KEYINPUT56), .C1(new_n809_), .C2(new_n800_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n817_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(new_n833_), .B2(new_n620_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n678_), .B1(new_n829_), .B2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n572_), .A2(new_n688_), .A3(new_n644_), .A4(new_n678_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(KEYINPUT117), .A3(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n623_), .A2(new_n572_), .A3(new_n644_), .A4(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT122), .B1(new_n836_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n833_), .A2(KEYINPUT57), .A3(new_n620_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n824_), .A2(new_n825_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n681_), .A3(new_n828_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(new_n846_), .C1(new_n818_), .C2(new_n830_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n842_), .B1(new_n847_), .B2(new_n586_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n789_), .B1(new_n843_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n490_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT123), .B(new_n855_), .C1(new_n836_), .C2(new_n842_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n851_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(KEYINPUT59), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n861_), .A2(new_n490_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n853_), .B1(new_n862_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g662(.A(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n572_), .B2(KEYINPUT60), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n851_), .B(new_n865_), .C1(KEYINPUT60), .C2(new_n864_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n861_), .A2(new_n643_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n864_), .ZN(G1341gat));
  AOI211_X1 g667(.A(KEYINPUT122), .B(new_n842_), .C1(new_n847_), .C2(new_n586_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n844_), .A2(new_n846_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n586_), .B1(new_n870_), .B2(new_n834_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n842_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n849_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n678_), .B(new_n788_), .C1(new_n869_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G127gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n857_), .A2(new_n858_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n586_), .A2(new_n875_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n879_), .B(new_n880_), .C1(new_n881_), .C2(new_n851_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n874_), .A2(KEYINPUT124), .A3(new_n875_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n878_), .A2(new_n882_), .A3(KEYINPUT125), .A4(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1342gat));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n860_), .B2(new_n640_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n892_), .B(new_n889_), .C1(new_n860_), .C2(new_n640_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n688_), .A2(new_n889_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n891_), .A2(new_n893_), .B1(new_n861_), .B2(new_n894_), .ZN(G1343gat));
  NAND2_X1  g694(.A1(new_n843_), .A2(new_n850_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n636_), .A2(new_n285_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n651_), .A2(new_n411_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(new_n206_), .A3(new_n490_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G141gat), .B1(new_n900_), .B2(new_n644_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1344gat));
  NAND3_X1  g703(.A1(new_n901_), .A2(new_n207_), .A3(new_n643_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G148gat), .B1(new_n900_), .B2(new_n572_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1345gat));
  XNOR2_X1  g706(.A(KEYINPUT61), .B(G155gat), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n900_), .A2(new_n586_), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n900_), .B2(new_n586_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1346gat));
  INV_X1    g710(.A(G162gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n900_), .A2(new_n912_), .A3(new_n682_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n901_), .A2(new_n641_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n912_), .B2(new_n914_), .ZN(G1347gat));
  AOI21_X1  g714(.A(new_n398_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n636_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n420_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n919_));
  OR3_X1    g718(.A1(new_n919_), .A2(KEYINPUT127), .A3(new_n644_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT127), .B1(new_n919_), .B2(new_n644_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n920_), .A2(G169gat), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n923_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n919_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n311_), .A3(new_n490_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(new_n925_), .A3(new_n927_), .ZN(G1348gat));
  AOI21_X1  g727(.A(G176gat), .B1(new_n926_), .B2(new_n643_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n420_), .B1(new_n843_), .B2(new_n850_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n917_), .A2(new_n572_), .A3(new_n299_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1349gat));
  NOR3_X1   g731(.A1(new_n919_), .A2(new_n302_), .A3(new_n586_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n930_), .A2(new_n636_), .A3(new_n678_), .A4(new_n916_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n323_), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n919_), .B2(new_n688_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n641_), .A2(new_n301_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n919_), .B2(new_n937_), .ZN(G1351gat));
  NAND3_X1  g737(.A1(new_n896_), .A2(new_n897_), .A3(new_n916_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n644_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n239_), .ZN(G1352gat));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n572_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n236_), .ZN(G1353gat));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n939_), .A2(new_n586_), .A3(new_n944_), .A4(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n898_), .A2(new_n678_), .A3(new_n916_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n944_), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n939_), .B2(new_n688_), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n640_), .A2(G218gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n939_), .B2(new_n950_), .ZN(G1355gat));
endmodule


