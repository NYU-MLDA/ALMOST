//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n938_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  INV_X1    g002(.A(G113gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT86), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G113gat), .ZN(new_n207_));
  INV_X1    g006(.A(G120gat), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n205_), .A2(new_n207_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G120gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n203_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n220_), .A2(new_n221_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n222_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(new_n218_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(KEYINPUT1), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT88), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n227_), .A2(KEYINPUT1), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n235_), .A2(new_n237_), .A3(new_n230_), .A4(new_n238_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n228_), .A2(new_n230_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n217_), .B1(new_n240_), .B2(KEYINPUT96), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n226_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n242_));
  AND4_X1   g041(.A1(new_n237_), .A2(new_n235_), .A3(new_n230_), .A4(new_n238_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n232_), .ZN(new_n244_));
  OAI211_X1 g043(.A(KEYINPUT96), .B(new_n242_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n211_), .A2(new_n216_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT4), .B1(new_n241_), .B2(new_n247_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n240_), .A2(KEYINPUT4), .A3(new_n246_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n202_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n202_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n241_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G85gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n251_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n240_), .A2(KEYINPUT96), .A3(new_n217_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n245_), .A2(new_n246_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n252_), .B1(new_n263_), .B2(new_n249_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n253_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n257_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OR3_X1    g065(.A1(new_n259_), .A2(new_n266_), .A3(KEYINPUT98), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT98), .B1(new_n259_), .B2(new_n266_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G43gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT31), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  OR2_X1    g074(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n276_));
  NAND2_X1  g075(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(G183gat), .B2(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n274_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT85), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT22), .ZN(new_n283_));
  AOI21_X1  g082(.A(G176gat), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G169gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT22), .B(G169gat), .ZN(new_n287_));
  INV_X1    g086(.A(G176gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT85), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n288_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT81), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT26), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT81), .B1(new_n299_), .B2(new_n303_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n301_), .A2(new_n304_), .A3(KEYINPUT82), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n295_), .A2(new_n296_), .B1(new_n299_), .B2(KEYINPUT81), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n302_), .A2(KEYINPUT26), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n298_), .A2(G190gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n306_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n294_), .B1(new_n305_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n275_), .A2(KEYINPUT23), .ZN(new_n315_));
  AND2_X1   g114(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n315_), .B1(new_n318_), .B2(new_n275_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n314_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n276_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n275_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n279_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n320_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT84), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n290_), .B1(new_n313_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT30), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n246_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n281_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT84), .B1(new_n325_), .B2(new_n326_), .ZN(new_n333_));
  AOI211_X1 g132(.A(new_n314_), .B(new_n320_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT82), .B1(new_n301_), .B2(new_n304_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n307_), .A2(new_n311_), .A3(new_n306_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n293_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT30), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n217_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n272_), .B1(new_n331_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  NAND3_X1  g145(.A1(new_n331_), .A2(new_n341_), .A3(new_n272_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n342_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G78gat), .B(G106gat), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n356_), .B(new_n242_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G22gat), .B(G50gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT28), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT92), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n355_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n355_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G204gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G197gat), .ZN(new_n369_));
  INV_X1    g168(.A(G197gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G204gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n371_), .A3(KEYINPUT90), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(KEYINPUT89), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G197gat), .B(G204gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT89), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(KEYINPUT90), .A4(KEYINPUT21), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n375_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n240_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(KEYINPUT29), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G228gat), .A2(G233gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT91), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n360_), .A2(KEYINPUT92), .A3(new_n361_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n385_), .A2(KEYINPUT91), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n384_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n367_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n366_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n392_), .A2(new_n364_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT93), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n280_), .B1(new_n398_), .B2(new_n323_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n399_), .B2(new_n320_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n309_), .A2(new_n310_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n293_), .B1(new_n401_), .B2(new_n297_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n326_), .B(KEYINPUT93), .C1(new_n278_), .C2(new_n280_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n283_), .A2(new_n285_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n405_), .A2(KEYINPUT94), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT94), .B1(new_n405_), .B2(new_n406_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n288_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n325_), .A2(new_n274_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n292_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n382_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n290_), .B(new_n382_), .C1(new_n313_), .C2(new_n328_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT20), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT19), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n404_), .A2(new_n382_), .A3(new_n411_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT95), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n329_), .A2(new_n413_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n404_), .A2(new_n382_), .A3(KEYINPUT95), .A4(new_n411_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT20), .A4(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT18), .B(G64gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G92gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G8gat), .B(G36gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  NAND3_X1  g228(.A1(new_n419_), .A2(new_n425_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n339_), .B2(new_n382_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n418_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n414_), .ZN(new_n434_));
  OAI211_X1 g233(.A(KEYINPUT20), .B(new_n420_), .C1(new_n339_), .C2(new_n382_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n418_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT27), .B(new_n430_), .C1(new_n437_), .C2(new_n429_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n429_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT20), .B(new_n424_), .C1(new_n339_), .C2(new_n382_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n420_), .A2(new_n421_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n433_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n433_), .B1(new_n432_), .B2(new_n414_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n439_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n430_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT27), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT99), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT99), .ZN(new_n449_));
  AOI211_X1 g248(.A(new_n449_), .B(KEYINPUT27), .C1(new_n445_), .C2(new_n430_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n396_), .B(new_n438_), .C1(new_n448_), .C2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(KEYINPUT100), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT100), .ZN(new_n453_));
  INV_X1    g252(.A(new_n438_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n419_), .A2(new_n425_), .A3(new_n429_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n429_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n447_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n449_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n446_), .A2(KEYINPUT99), .A3(new_n447_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n454_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n453_), .B1(new_n460_), .B2(new_n396_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n269_), .B(new_n353_), .C1(new_n452_), .C2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n429_), .A2(KEYINPUT32), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n419_), .A2(new_n425_), .A3(new_n463_), .ZN(new_n464_));
  OAI221_X1 g263(.A(new_n464_), .B1(new_n437_), .B2(new_n463_), .C1(new_n259_), .C2(new_n266_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n455_), .A2(new_n456_), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT33), .B(new_n258_), .C1(new_n251_), .C2(new_n253_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT97), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT97), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n266_), .A2(new_n469_), .A3(KEYINPUT33), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n258_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n466_), .A2(new_n468_), .A3(new_n470_), .A4(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n263_), .A2(new_n252_), .A3(new_n249_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n202_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n258_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n465_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n396_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n396_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n460_), .A2(new_n269_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n348_), .A2(new_n351_), .A3(KEYINPUT87), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT87), .B1(new_n348_), .B2(new_n351_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n462_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT74), .B(G29gat), .ZN(new_n489_));
  INV_X1    g288(.A(G36gat), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n490_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n488_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(KEYINPUT15), .A3(new_n494_), .ZN(new_n499_));
  INV_X1    g298(.A(G1gat), .ZN(new_n500_));
  INV_X1    g299(.A(G8gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT77), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT77), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G1gat), .B(G8gat), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n503_), .A2(new_n507_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n497_), .A2(new_n499_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n498_), .A2(new_n494_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n510_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT78), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR4_X1   g316(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G141gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT79), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(new_n204_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n511_), .A2(new_n517_), .A3(new_n514_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n498_), .A2(new_n494_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n517_), .B1(new_n514_), .B2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n526_), .A2(KEYINPUT78), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n519_), .B(new_n523_), .C1(new_n524_), .C2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n523_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n511_), .A2(new_n514_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n530_), .A2(new_n516_), .B1(new_n526_), .B2(KEYINPUT78), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n531_), .B2(new_n518_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n528_), .A2(KEYINPUT80), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT80), .B1(new_n528_), .B2(new_n532_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G71gat), .ZN(new_n536_));
  INV_X1    g335(.A(G78gat), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n537_), .A2(KEYINPUT69), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(KEYINPUT69), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT69), .B(G78gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(G71gat), .ZN(new_n542_));
  OR2_X1    g341(.A1(G57gat), .A2(G64gat), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G57gat), .A2(G64gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n540_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT70), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n544_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT70), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n540_), .A2(new_n542_), .A3(new_n550_), .A4(new_n546_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n549_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(G99gat), .ZN(new_n555_));
  INV_X1    g354(.A(G106gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT67), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n558_), .B1(G99gat), .B2(G106gat), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT7), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT68), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT68), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n557_), .A2(new_n559_), .A3(new_n563_), .A4(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT6), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT66), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n562_), .A2(new_n564_), .A3(new_n566_), .A4(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G85gat), .B(G92gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n572_), .A2(KEYINPUT8), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT8), .B1(new_n572_), .B2(new_n574_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(G85gat), .A3(G92gat), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n566_), .B(new_n579_), .C1(new_n578_), .C2(new_n573_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT65), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT10), .B(G99gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n583_), .B2(new_n556_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n582_), .A2(KEYINPUT65), .A3(G106gat), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n580_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT71), .B1(new_n577_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n572_), .A2(new_n574_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT8), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n572_), .A2(KEYINPUT8), .A3(new_n574_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n590_), .A2(KEYINPUT71), .A3(new_n591_), .A4(new_n586_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(KEYINPUT12), .B(new_n554_), .C1(new_n587_), .C2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n591_), .A3(new_n586_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT12), .B1(new_n595_), .B2(new_n554_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n554_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G230gat), .A2(G233gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT64), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n594_), .A2(new_n598_), .A3(KEYINPUT72), .A4(new_n600_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n600_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(new_n554_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(new_n597_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n603_), .A2(new_n604_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n368_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n288_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n609_), .A2(new_n613_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT13), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n614_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n535_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n497_), .A2(new_n499_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n587_), .B2(new_n593_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT73), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT34), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT35), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT76), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n495_), .A2(new_n496_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n590_), .A2(new_n630_), .A3(new_n591_), .A4(new_n586_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n626_), .A2(KEYINPUT35), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(KEYINPUT76), .A3(KEYINPUT35), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n623_), .A2(new_n629_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n629_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n622_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT71), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n595_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n640_), .B2(new_n592_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n641_), .B2(new_n634_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(G134gat), .ZN(new_n644_));
  INV_X1    g443(.A(G162gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n636_), .A2(new_n642_), .A3(KEYINPUT36), .A4(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(KEYINPUT36), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n636_), .A2(new_n642_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT75), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT75), .B(new_n649_), .C1(new_n636_), .C2(new_n642_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n648_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT37), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT37), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n657_), .B(new_n648_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(G231gat), .A2(G233gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n513_), .B(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(new_n554_), .Z(new_n662_));
  INV_X1    g461(.A(KEYINPUT17), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G183gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(G211gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(G127gat), .B(G155gat), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n665_), .B(new_n666_), .Z(new_n667_));
  NOR3_X1   g466(.A1(new_n662_), .A2(new_n663_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(KEYINPUT17), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n662_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n659_), .A2(new_n671_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n487_), .A2(new_n621_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n269_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n500_), .A3(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT38), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n655_), .A2(new_n671_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n487_), .A2(new_n677_), .A3(new_n621_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G1gat), .B1(new_n678_), .B2(new_n269_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1324gat));
  OAI21_X1  g479(.A(G8gat), .B1(new_n678_), .B2(new_n460_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT101), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n683_), .B(G8gat), .C1(new_n678_), .C2(new_n460_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(KEYINPUT39), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n460_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n673_), .A2(new_n501_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n681_), .A2(KEYINPUT101), .A3(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n687_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT102), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n685_), .A2(new_n692_), .A3(new_n687_), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n691_), .A2(KEYINPUT40), .A3(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1325gat));
  OAI21_X1  g497(.A(G15gat), .B1(new_n678_), .B2(new_n485_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT103), .Z(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT41), .ZN(new_n701_));
  INV_X1    g500(.A(G15gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n485_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n673_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1326gat));
  OAI21_X1  g504(.A(G22gat), .B1(new_n678_), .B2(new_n396_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT42), .ZN(new_n707_));
  INV_X1    g506(.A(G22gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n673_), .A2(new_n708_), .A3(new_n480_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1327gat));
  NAND2_X1  g509(.A1(new_n655_), .A2(new_n671_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n487_), .A2(new_n621_), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n487_), .A2(KEYINPUT105), .A3(new_n621_), .A4(new_n712_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G29gat), .B1(new_n717_), .B2(new_n674_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n656_), .A2(KEYINPUT104), .A3(new_n658_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT104), .B1(new_n656_), .B2(new_n658_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n719_), .B1(new_n487_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n451_), .A2(KEYINPUT100), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n460_), .A2(new_n453_), .A3(new_n396_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n674_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n726_), .A2(new_n353_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n659_), .A2(new_n719_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n671_), .B(new_n621_), .C1(new_n723_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n659_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n656_), .A2(KEYINPUT104), .A3(new_n658_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n727_), .B2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n487_), .A2(new_n659_), .A3(new_n719_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(KEYINPUT44), .A3(new_n671_), .A4(new_n621_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n732_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(G29gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n718_), .B1(new_n742_), .B2(new_n674_), .ZN(G1328gat));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n715_), .A2(new_n490_), .A3(new_n686_), .A4(new_n716_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT106), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(KEYINPUT106), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n748_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(KEYINPUT45), .A3(new_n746_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n732_), .A2(new_n740_), .A3(new_n686_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G36gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT107), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT108), .Z(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n749_), .A2(new_n751_), .A3(new_n757_), .A4(new_n753_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1329gat));
  INV_X1    g560(.A(G43gat), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n352_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n732_), .A2(new_n740_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT109), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n732_), .A2(new_n740_), .A3(new_n766_), .A4(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n717_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n762_), .B1(new_n769_), .B2(new_n485_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n772_), .A3(new_n770_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1330gat));
  AOI21_X1  g575(.A(G50gat), .B1(new_n717_), .B2(new_n480_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n480_), .A2(G50gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n741_), .B2(new_n778_), .ZN(G1331gat));
  NAND2_X1  g578(.A1(new_n617_), .A2(new_n620_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n535_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(new_n487_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n672_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G57gat), .B1(new_n784_), .B2(new_n674_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n783_), .A2(new_n677_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(G57gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n674_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT111), .ZN(G1332gat));
  INV_X1    g588(.A(G64gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n786_), .B2(new_n686_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT48), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n784_), .A2(new_n790_), .A3(new_n686_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1333gat));
  NAND3_X1  g593(.A1(new_n784_), .A2(new_n536_), .A3(new_n703_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n786_), .A2(new_n703_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G71gat), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n797_), .A2(KEYINPUT112), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(KEYINPUT112), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(KEYINPUT49), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT49), .B1(new_n798_), .B2(new_n799_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n795_), .B1(new_n800_), .B2(new_n801_), .ZN(G1334gat));
  AOI21_X1  g601(.A(new_n537_), .B1(new_n786_), .B2(new_n480_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT50), .Z(new_n804_));
  NAND3_X1  g603(.A1(new_n784_), .A2(new_n537_), .A3(new_n480_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1335gat));
  AND2_X1   g605(.A1(new_n783_), .A2(new_n712_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G85gat), .B1(new_n807_), .B2(new_n674_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n670_), .B1(new_n739_), .B2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n782_), .C1(new_n809_), .C2(new_n739_), .ZN(new_n811_));
  INV_X1    g610(.A(G85gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n808_), .B1(new_n813_), .B2(new_n674_), .ZN(G1336gat));
  AOI21_X1  g613(.A(G92gat), .B1(new_n807_), .B2(new_n686_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n811_), .A2(new_n460_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g616(.A(G99gat), .B1(new_n811_), .B2(new_n485_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n807_), .A2(new_n583_), .A3(new_n353_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT114), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT115), .A3(KEYINPUT51), .ZN(new_n822_));
  NAND2_X1  g621(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1338gat));
  NAND3_X1  g624(.A1(new_n807_), .A2(new_n556_), .A3(new_n480_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n739_), .A2(new_n671_), .A3(new_n480_), .A4(new_n782_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G106gat), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n828_), .A2(KEYINPUT52), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(KEYINPUT52), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n826_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT53), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(new_n826_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1339gat));
  OAI211_X1 g634(.A(new_n674_), .B(new_n353_), .C1(new_n452_), .C2(new_n461_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT118), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n613_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT55), .B1(new_n603_), .B2(new_n604_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n594_), .A2(new_n598_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n605_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n601_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n839_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n839_), .B(new_n846_), .C1(new_n840_), .C2(new_n844_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n848_), .A2(new_n781_), .A3(new_n614_), .A4(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n528_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n516_), .B1(new_n514_), .B2(new_n525_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n523_), .B1(new_n530_), .B2(new_n517_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n850_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n655_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n859_), .B(new_n655_), .C1(new_n850_), .C2(new_n855_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n845_), .A2(KEYINPUT56), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n614_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n854_), .B1(new_n845_), .B2(KEYINPUT56), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT58), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n862_), .B(new_n868_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n659_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n670_), .B1(new_n861_), .B2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n672_), .A2(new_n535_), .A3(new_n780_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT54), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n672_), .A2(new_n780_), .A3(new_n874_), .A4(new_n535_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n838_), .B1(new_n871_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n838_), .B(new_n881_), .C1(new_n871_), .C2(new_n877_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n879_), .A2(G113gat), .A3(new_n781_), .A4(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n204_), .B1(new_n878_), .B2(new_n535_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1340gat));
  INV_X1    g684(.A(new_n878_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n208_), .B1(new_n780_), .B2(KEYINPUT60), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n886_), .B(new_n887_), .C1(KEYINPUT60), .C2(new_n208_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n780_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n879_), .A2(new_n889_), .A3(new_n882_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n890_), .B2(new_n208_), .ZN(G1341gat));
  INV_X1    g690(.A(G127gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n878_), .B2(new_n671_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n893_), .A2(KEYINPUT120), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(KEYINPUT120), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n879_), .A2(G127gat), .A3(new_n670_), .A4(new_n882_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(G1342gat));
  AOI21_X1  g696(.A(G134gat), .B1(new_n886_), .B2(new_n655_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n879_), .A2(new_n882_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n659_), .A2(G134gat), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT121), .Z(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n899_), .B2(new_n901_), .ZN(G1343gat));
  OAI211_X1 g701(.A(new_n674_), .B(new_n460_), .C1(new_n871_), .C2(new_n877_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n703_), .A2(new_n396_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n781_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n889_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n670_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  NAND2_X1  g712(.A1(new_n861_), .A2(new_n870_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n671_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n269_), .B1(new_n915_), .B2(new_n876_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n736_), .A2(new_n645_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n916_), .A2(new_n460_), .A3(new_n904_), .A4(new_n917_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n903_), .A2(new_n857_), .A3(new_n905_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(G162gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT122), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n918_), .B(new_n922_), .C1(new_n919_), .C2(G162gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n485_), .A2(new_n674_), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n686_), .B(new_n925_), .C1(new_n871_), .C2(new_n877_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n480_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n927_), .B(new_n781_), .C1(new_n408_), .C2(new_n407_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n925_), .A2(new_n781_), .A3(new_n686_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT123), .Z(new_n930_));
  OAI211_X1 g729(.A(new_n396_), .B(new_n930_), .C1(new_n871_), .C2(new_n877_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n931_), .A2(new_n932_), .A3(G169gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n931_), .B2(G169gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n928_), .B1(new_n933_), .B2(new_n934_), .ZN(G1348gat));
  NAND2_X1  g734(.A1(new_n927_), .A2(new_n889_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g736(.A1(new_n926_), .A2(new_n671_), .A3(new_n480_), .ZN(new_n938_));
  MUX2_X1   g737(.A(G183gat), .B(new_n297_), .S(new_n938_), .Z(G1350gat));
  AOI21_X1  g738(.A(new_n460_), .B1(new_n915_), .B2(new_n876_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n655_), .A2(new_n401_), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n940_), .A2(new_n396_), .A3(new_n925_), .A4(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n659_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n926_), .A2(new_n480_), .A3(new_n943_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n942_), .B1(new_n944_), .B2(new_n302_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(KEYINPUT124), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n942_), .B(new_n947_), .C1(new_n944_), .C2(new_n302_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(G1351gat));
  NAND2_X1  g748(.A1(new_n904_), .A2(new_n269_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n940_), .A2(new_n951_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n952_), .A2(new_n535_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(new_n370_), .ZN(G1352gat));
  OAI22_X1  g753(.A1(new_n952_), .A2(new_n780_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n955_));
  NAND2_X1  g754(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n956_), .B(KEYINPUT126), .Z(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n955_), .A2(new_n958_), .ZN(new_n959_));
  OAI221_X1 g758(.A(new_n957_), .B1(KEYINPUT125), .B2(G204gat), .C1(new_n952_), .C2(new_n780_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(G1353gat));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  NAND4_X1  g763(.A1(new_n940_), .A2(new_n670_), .A3(new_n951_), .A4(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n962_), .B1(new_n965_), .B2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n686_), .B1(new_n871_), .B2(new_n877_), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n969_), .A2(new_n671_), .A3(new_n950_), .ZN(new_n970_));
  NAND4_X1  g769(.A1(new_n970_), .A2(KEYINPUT127), .A3(new_n964_), .A4(new_n966_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n963_), .B1(new_n952_), .B2(new_n671_), .ZN(new_n972_));
  AND3_X1   g771(.A1(new_n968_), .A2(new_n971_), .A3(new_n972_), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974_));
  NOR3_X1   g773(.A1(new_n952_), .A2(new_n974_), .A3(new_n943_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n940_), .A2(new_n655_), .A3(new_n951_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n975_), .B1(new_n974_), .B2(new_n976_), .ZN(G1355gat));
endmodule


