//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  XOR2_X1   g000(.A(G22gat), .B(G50gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G155gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT84), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G155gat), .B2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n204_), .B2(new_n205_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G155gat), .A3(G162gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G141gat), .B(G148gat), .Z(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI22_X1  g016(.A1(KEYINPUT85), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n217_), .A2(new_n218_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n206_), .A2(new_n208_), .B1(G155gat), .B2(G162gat), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n213_), .A2(new_n214_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n227_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n203_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n227_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n206_), .A2(new_n208_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n210_), .A2(new_n212_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n214_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n223_), .A2(new_n224_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n232_), .B1(new_n237_), .B2(KEYINPUT29), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(new_n202_), .A3(new_n228_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G197gat), .B(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G218gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G211gat), .ZN(new_n245_));
  INV_X1    g044(.A(G211gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G218gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT88), .ZN(new_n250_));
  INV_X1    g049(.A(G204gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(G197gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT21), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(KEYINPUT88), .B2(new_n241_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(G197gat), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G204gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n245_), .B(new_n247_), .C1(new_n258_), .C2(KEYINPUT21), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n249_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(G228gat), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n260_), .B(new_n264_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT90), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n267_));
  OAI21_X1  g066(.A(new_n260_), .B1(new_n225_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n264_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n267_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n248_), .B1(new_n242_), .B2(new_n241_), .ZN(new_n272_));
  OAI211_X1 g071(.A(KEYINPUT21), .B(new_n252_), .C1(new_n258_), .C2(new_n250_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n272_), .A2(new_n273_), .B1(new_n248_), .B2(new_n243_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n266_), .B(new_n269_), .C1(new_n271_), .C2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n265_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G78gat), .B(G106gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n240_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(new_n265_), .C1(new_n270_), .C2(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT92), .ZN(new_n282_));
  INV_X1    g081(.A(new_n265_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n269_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT90), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n285_), .B2(new_n275_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n280_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n240_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n277_), .A2(new_n278_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(new_n281_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n289_), .B1(new_n292_), .B2(KEYINPUT91), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  AOI211_X1 g093(.A(new_n294_), .B(new_n290_), .C1(new_n291_), .C2(new_n281_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT93), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n281_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n286_), .A2(new_n280_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n240_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n294_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n292_), .A2(KEYINPUT91), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT93), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .A4(new_n289_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G15gat), .B(G43gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT81), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G227gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT82), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G71gat), .B(G99gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(KEYINPUT76), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n314_), .B2(KEYINPUT23), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT25), .B(G183gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G190gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n319_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(KEYINPUT77), .A2(G176gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT22), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT22), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G169gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(KEYINPUT77), .A2(G176gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n334_), .A2(new_n336_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n339_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(new_n333_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G169gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT78), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n324_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n315_), .A2(new_n313_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT79), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352_));
  AOI211_X1 g151(.A(new_n352_), .B(new_n349_), .C1(new_n315_), .C2(new_n313_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n332_), .B1(new_n347_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n357_), .A2(new_n358_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n311_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n359_), .B2(new_n311_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n363_), .A2(new_n364_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT31), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n362_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  AND4_X1   g170(.A1(new_n371_), .A2(new_n367_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n367_), .B1(new_n225_), .B2(new_n371_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT4), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n237_), .A2(new_n375_), .A3(new_n367_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n370_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n370_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n372_), .A2(new_n373_), .A3(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G85gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT0), .B(G57gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  OR3_X1    g182(.A1(new_n377_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n383_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n319_), .A2(new_n350_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n324_), .A2(new_n340_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n326_), .A2(new_n320_), .B1(new_n315_), .B2(new_n313_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n389_), .A2(new_n390_), .B1(new_n331_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n392_), .B2(new_n274_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n355_), .A2(new_n260_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT19), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT94), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n274_), .B(new_n332_), .C1(new_n347_), .C2(new_n354_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(KEYINPUT20), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n392_), .A2(new_n274_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n399_), .A3(KEYINPUT20), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n398_), .B1(new_n405_), .B2(new_n396_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G8gat), .B(G36gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n387_), .B1(new_n406_), .B2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n405_), .A2(new_n396_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n397_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n411_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n404_), .A2(new_n403_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n396_), .B1(new_n418_), .B2(new_n401_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n398_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n419_), .A2(new_n412_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n412_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n417_), .B1(KEYINPUT27), .B2(new_n423_), .ZN(new_n424_));
  NOR4_X1   g223(.A1(new_n304_), .A2(new_n369_), .A3(new_n386_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT97), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n385_), .B2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT33), .B(new_n383_), .C1(new_n377_), .C2(new_n379_), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n237_), .A2(KEYINPUT96), .B1(new_n365_), .B2(new_n366_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n225_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n370_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT98), .B1(new_n432_), .B2(new_n383_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n378_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n383_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT98), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n374_), .A2(new_n370_), .A3(new_n376_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n433_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n429_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n428_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n385_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n423_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n406_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n414_), .A2(new_n415_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n386_), .B(new_n445_), .C1(new_n446_), .C2(new_n444_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n296_), .A2(new_n443_), .A3(new_n303_), .A4(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n369_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n422_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n406_), .A2(new_n412_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n452_), .A2(new_n387_), .B1(new_n416_), .B2(new_n413_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n386_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n453_), .A2(new_n454_), .B1(new_n296_), .B2(new_n303_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT99), .B1(new_n449_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n304_), .B1(new_n386_), .B2(new_n424_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n448_), .A4(new_n369_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n425_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G29gat), .B(G36gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT68), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G43gat), .B(G50gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT69), .B(G15gat), .ZN(new_n465_));
  INV_X1    g264(.A(G22gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT14), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT70), .B(G8gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(G1gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G8gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n473_), .A2(new_n475_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n464_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n473_), .A2(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n473_), .A2(new_n475_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n464_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n473_), .B(new_n474_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n464_), .B(KEYINPUT15), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n484_), .B(KEYINPUT74), .Z(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n478_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G169gat), .B(G197gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n486_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n460_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G106gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT10), .B(G99gat), .Z(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n508_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n507_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT65), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n510_), .A2(new_n511_), .ZN(new_n518_));
  INV_X1    g317(.A(G99gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n505_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT66), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n520_), .B(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n518_), .B1(new_n523_), .B2(new_n504_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT8), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n488_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  OAI221_X1 g329(.A(new_n527_), .B1(KEYINPUT35), .B2(new_n530_), .C1(new_n481_), .C2(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(KEYINPUT35), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G190gat), .B(G218gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT36), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n533_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n534_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n537_), .B(KEYINPUT36), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT37), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n539_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n541_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n534_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n544_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT16), .ZN(new_n552_));
  XOR2_X1   g351(.A(G183gat), .B(G211gat), .Z(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT72), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n487_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n562_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n556_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n558_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n558_), .B2(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n554_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n570_), .A2(new_n571_), .A3(KEYINPUT73), .ZN(new_n575_));
  INV_X1    g374(.A(new_n554_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n579_), .B(new_n572_), .C1(new_n574_), .C2(new_n577_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n550_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n526_), .A2(new_n568_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n517_), .A2(new_n567_), .A3(new_n525_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT12), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT12), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n526_), .A2(new_n587_), .A3(new_n568_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n583_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G120gat), .B(G148gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT5), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  OR3_X1    g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(KEYINPUT13), .A3(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n581_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n501_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(G1gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n386_), .B(KEYINPUT100), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT102), .B1(new_n540_), .B2(new_n543_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n546_), .A2(new_n611_), .A3(new_n548_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n460_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n601_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(KEYINPUT101), .A3(new_n499_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n578_), .A2(new_n580_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n601_), .B2(new_n500_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n617_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n615_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n454_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n607_), .A2(new_n608_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n609_), .A2(new_n624_), .A3(new_n625_), .ZN(G1324gat));
  OAI21_X1  g425(.A(G8gat), .B1(new_n623_), .B2(new_n453_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT39), .ZN(new_n628_));
  INV_X1    g427(.A(new_n469_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n603_), .A2(new_n424_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT103), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n603_), .A2(new_n632_), .A3(new_n424_), .A4(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n628_), .B2(new_n634_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(new_n369_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n615_), .A2(new_n622_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G15gat), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT105), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT105), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT41), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT41), .ZN(new_n646_));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n603_), .A2(new_n647_), .A3(new_n639_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT106), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n646_), .A3(new_n649_), .ZN(G1326gat));
  XNOR2_X1  g449(.A(new_n304_), .B(KEYINPUT107), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n603_), .A2(new_n466_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G22gat), .B1(new_n623_), .B2(new_n651_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n456_), .A2(new_n459_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n425_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  INV_X1    g460(.A(new_n550_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n550_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n617_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT44), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  AOI211_X1 g468(.A(new_n669_), .B(new_n666_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n605_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n614_), .A2(new_n618_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n601_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n501_), .A2(new_n386_), .A3(new_n675_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n671_), .A2(new_n673_), .B1(new_n676_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n671_), .B2(new_n424_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n453_), .A2(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n501_), .A2(new_n675_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT108), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n501_), .A2(new_n684_), .A3(new_n675_), .A4(new_n681_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT45), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(KEYINPUT45), .A3(new_n685_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n678_), .B1(new_n680_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n688_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n686_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n668_), .A2(new_n670_), .A3(new_n453_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n692_), .B(KEYINPUT46), .C1(new_n693_), .C2(new_n679_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(G43gat), .ZN(new_n696_));
  NOR4_X1   g495(.A1(new_n668_), .A2(new_n670_), .A3(new_n696_), .A4(new_n369_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n501_), .A2(new_n675_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n698_), .B2(new_n369_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT47), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n671_), .A2(G43gat), .A3(new_n639_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n699_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1330gat));
  INV_X1    g504(.A(new_n304_), .ZN(new_n706_));
  INV_X1    g505(.A(G50gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n501_), .A2(new_n652_), .A3(new_n675_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n671_), .A2(new_n708_), .B1(new_n709_), .B2(new_n707_), .ZN(G1331gat));
  NAND2_X1  g509(.A1(new_n601_), .A2(new_n500_), .ZN(new_n711_));
  NOR4_X1   g510(.A1(new_n460_), .A2(new_n618_), .A3(new_n614_), .A4(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(G57gat), .A3(new_n386_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n714_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n460_), .A2(new_n499_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n581_), .A2(new_n616_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n606_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n715_), .A2(new_n716_), .A3(new_n721_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n712_), .B2(new_n424_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT48), .Z(new_n725_));
  NAND2_X1  g524(.A1(new_n424_), .A2(new_n723_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT110), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n719_), .B2(new_n727_), .ZN(G1333gat));
  INV_X1    g527(.A(G71gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n712_), .B2(new_n639_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT49), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n639_), .A2(new_n729_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT111), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n719_), .B2(new_n733_), .ZN(G1334gat));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n712_), .B2(new_n652_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT50), .Z(new_n737_));
  NAND3_X1  g536(.A1(new_n720_), .A2(new_n735_), .A3(new_n652_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n619_), .A2(new_n711_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n661_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n460_), .A2(KEYINPUT43), .A3(new_n550_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n665_), .A2(KEYINPUT113), .A3(new_n740_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n386_), .A2(G85gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT114), .ZN(new_n749_));
  NOR4_X1   g548(.A1(new_n460_), .A2(new_n674_), .A3(new_n499_), .A4(new_n616_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n606_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT112), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT112), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n747_), .A2(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  INV_X1    g553(.A(G92gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n755_), .A3(new_n424_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n453_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n755_), .ZN(G1337gat));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n639_), .A2(new_n506_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n750_), .B2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n369_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n519_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n761_), .C1(new_n762_), .C2(new_n519_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n750_), .A2(new_n505_), .A3(new_n304_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n665_), .A2(new_n304_), .A3(new_n740_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n768_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  NOR2_X1   g576(.A1(new_n424_), .A2(new_n605_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(new_n369_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n483_), .A2(new_n490_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n490_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n489_), .A2(new_n478_), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n496_), .A3(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n498_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n597_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n597_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n499_), .A2(new_n595_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n589_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n586_), .A2(new_n583_), .A3(new_n588_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n594_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n589_), .B2(new_n792_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n797_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n791_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n613_), .B1(new_n790_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n785_), .A2(new_n595_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n800_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n798_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n550_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n804_), .B(KEYINPUT58), .C1(new_n805_), .C2(new_n798_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n802_), .A2(new_n803_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT57), .B(new_n613_), .C1(new_n790_), .C2(new_n801_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n619_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n602_), .A2(new_n500_), .A3(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n581_), .A2(new_n499_), .A3(new_n601_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n813_), .B(new_n814_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n706_), .B(new_n780_), .C1(new_n812_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(KEYINPUT59), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n817_), .A2(new_n818_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n815_), .ZN(new_n824_));
  NOR4_X1   g623(.A1(new_n581_), .A2(new_n601_), .A3(new_n499_), .A4(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n802_), .A2(new_n803_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n808_), .A2(new_n809_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n811_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n618_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n706_), .A3(new_n780_), .A4(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n500_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n822_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n820_), .B2(new_n500_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT119), .B(new_n834_), .C1(new_n820_), .C2(new_n500_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n836_), .A2(new_n839_), .A3(new_n840_), .ZN(G1340gat));
  NAND3_X1  g640(.A1(new_n822_), .A2(new_n601_), .A3(new_n833_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G120gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n820_), .ZN(new_n844_));
  INV_X1    g643(.A(G120gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n616_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(new_n846_), .C1(KEYINPUT60), .C2(new_n845_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n847_), .ZN(G1341gat));
  NAND3_X1  g647(.A1(new_n822_), .A2(new_n619_), .A3(new_n833_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G127gat), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n820_), .A2(G127gat), .A3(new_n618_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n550_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n822_), .A2(new_n833_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n820_), .B2(new_n613_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT121), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n858_), .B(new_n853_), .C1(new_n820_), .C2(new_n613_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n855_), .A2(new_n857_), .A3(new_n859_), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n706_), .A2(new_n639_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n778_), .B(new_n861_), .C1(new_n812_), .C2(new_n819_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n500_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n616_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(G148gat), .Z(G1345gat));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n862_), .B2(new_n618_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n861_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n870_), .A2(KEYINPUT122), .A3(new_n619_), .A4(new_n778_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n868_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1346gat));
  NOR3_X1   g674(.A1(new_n862_), .A2(new_n205_), .A3(new_n550_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n205_), .B1(new_n862_), .B2(new_n613_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT123), .B(new_n205_), .C1(new_n862_), .C2(new_n613_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(G1347gat));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n369_), .A2(new_n606_), .A3(new_n453_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n652_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n499_), .B(new_n885_), .C1(new_n812_), .C2(new_n819_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n886_), .B2(G169gat), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n888_));
  INV_X1    g687(.A(new_n886_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n887_), .A2(new_n888_), .B1(new_n345_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(G169gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT125), .ZN(new_n892_));
  INV_X1    g691(.A(new_n888_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n891_), .A2(KEYINPUT125), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n890_), .B1(new_n894_), .B2(new_n895_), .ZN(G1348gat));
  NAND2_X1  g695(.A1(new_n831_), .A2(new_n885_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n601_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n304_), .B(new_n884_), .C1(new_n826_), .C2(new_n830_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n601_), .A2(G176gat), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n899_), .A2(new_n344_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  AOI21_X1  g701(.A(G183gat), .B1(new_n900_), .B2(new_n619_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n897_), .A2(new_n329_), .A3(new_n618_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n897_), .B2(new_n550_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n614_), .A2(new_n330_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n897_), .B2(new_n907_), .ZN(G1351gat));
  NOR2_X1   g707(.A1(new_n453_), .A2(new_n386_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n870_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n500_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n256_), .ZN(G1352gat));
  NOR2_X1   g711(.A1(new_n251_), .A2(KEYINPUT126), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n251_), .A2(KEYINPUT126), .ZN(new_n914_));
  OAI22_X1  g713(.A1(new_n910_), .A2(new_n616_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n910_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n601_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n917_), .B2(new_n913_), .ZN(G1353gat));
  XOR2_X1   g717(.A(KEYINPUT63), .B(G211gat), .Z(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n619_), .A3(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n910_), .B2(new_n618_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n910_), .B2(new_n550_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n614_), .A2(new_n244_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n910_), .B2(new_n925_), .ZN(G1355gat));
endmodule


