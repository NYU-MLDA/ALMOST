//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G71gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G99gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT25), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G190gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n211_), .A2(new_n213_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n209_), .A2(new_n218_), .A3(new_n222_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT22), .B1(new_n228_), .B2(new_n224_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n225_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n210_), .A2(new_n214_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n219_), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n206_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n227_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n205_), .B(new_n239_), .Z(new_n240_));
  INV_X1    g039(.A(G134gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G127gat), .ZN(new_n242_));
  INV_X1    g041(.A(G127gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G134gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G120gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G113gat), .ZN(new_n247_));
  INV_X1    g046(.A(G113gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G120gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT85), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n250_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n242_), .A2(new_n244_), .A3(new_n247_), .A4(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(new_n254_), .B2(KEYINPUT85), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n240_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G15gat), .B(G43gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT84), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT30), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT31), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n256_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G22gat), .B(G50gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT87), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT2), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271_));
  INV_X1    g070(.A(G141gat), .ZN(new_n272_));
  INV_X1    g071(.A(G148gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n266_), .A2(new_n269_), .A3(new_n270_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G155gat), .ZN(new_n276_));
  INV_X1    g075(.A(G162gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT86), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(G155gat), .B2(G162gat), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n278_), .A2(new_n280_), .B1(G155gat), .B2(G162gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT1), .B1(new_n276_), .B2(new_n277_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(G155gat), .A3(G162gat), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n279_), .A2(G155gat), .A3(G162gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT86), .B1(new_n276_), .B2(new_n277_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n282_), .B(new_n284_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G141gat), .B(G148gat), .Z(new_n288_));
  AOI22_X1  g087(.A1(new_n275_), .A2(new_n281_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n262_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n274_), .B(new_n270_), .C1(new_n268_), .C2(new_n267_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n269_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n281_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n278_), .A2(new_n280_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n282_), .A2(new_n284_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  AND4_X1   g096(.A1(new_n290_), .A2(new_n294_), .A3(new_n297_), .A4(new_n262_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n291_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n289_), .A2(new_n290_), .A3(new_n262_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n297_), .A3(new_n290_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n262_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n299_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT91), .B1(new_n301_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT92), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n290_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n312_));
  OAI211_X1 g111(.A(KEYINPUT21), .B(new_n310_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT21), .ZN(new_n314_));
  INV_X1    g113(.A(G218gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G211gat), .ZN(new_n316_));
  INV_X1    g115(.A(G211gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G218gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n314_), .B1(new_n319_), .B2(KEYINPUT89), .ZN(new_n320_));
  AND2_X1   g119(.A1(G197gat), .A2(G204gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G197gat), .A2(G204gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n311_), .B2(KEYINPUT21), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n313_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(G78gat), .B1(new_n309_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G106gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n310_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT21), .B1(new_n311_), .B2(new_n312_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n329_), .B1(new_n332_), .B2(new_n313_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n328_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G78gat), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n336_), .B(new_n325_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n325_), .A2(KEYINPUT90), .ZN(new_n338_));
  INV_X1    g137(.A(new_n334_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(G106gat), .A3(new_n339_), .ZN(new_n340_));
  AND4_X1   g139(.A1(new_n327_), .A2(new_n335_), .A3(new_n337_), .A4(new_n340_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n335_), .A2(new_n340_), .B1(new_n327_), .B2(new_n337_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n300_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n302_), .A2(new_n305_), .A3(new_n299_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT91), .A3(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n308_), .A2(new_n343_), .A3(new_n347_), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n335_), .A2(new_n340_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n327_), .A2(new_n337_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n335_), .A2(new_n327_), .A3(new_n337_), .A4(new_n340_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n347_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n349_), .B1(new_n348_), .B2(KEYINPUT91), .ZN(new_n357_));
  AOI211_X1 g156(.A(new_n345_), .B(KEYINPUT92), .C1(new_n344_), .C2(new_n346_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT20), .B1(new_n239_), .B2(new_n325_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT94), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n212_), .A2(G183gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n215_), .A2(new_n217_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT94), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n226_), .A2(new_n235_), .A3(new_n219_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n207_), .A2(new_n208_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT95), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n237_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G169gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n207_), .B1(new_n375_), .B2(new_n225_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT95), .A4(new_n219_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n372_), .A2(new_n378_), .B1(new_n332_), .B2(new_n313_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OR3_X1    g182(.A1(new_n361_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n239_), .B2(new_n325_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n372_), .A2(new_n378_), .A3(new_n332_), .A4(new_n313_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT102), .ZN(new_n391_));
  XOR2_X1   g190(.A(G8gat), .B(G36gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT18), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT32), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n390_), .A2(new_n391_), .A3(new_n397_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n361_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(new_n388_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT102), .B1(new_n400_), .B2(new_n396_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n383_), .B1(new_n361_), .B2(new_n379_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n386_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n396_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n398_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n294_), .A2(new_n297_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n255_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(KEYINPUT4), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT97), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n245_), .A2(new_n250_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n242_), .A2(new_n244_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT97), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n294_), .A3(new_n297_), .A4(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(KEYINPUT4), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT98), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT98), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n407_), .A2(new_n414_), .A3(new_n417_), .A4(KEYINPUT4), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT99), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n407_), .A2(new_n423_), .A3(new_n414_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G85gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT0), .B(G57gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n423_), .B(new_n408_), .C1(new_n416_), .C2(new_n418_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n424_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n405_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n402_), .A2(new_n395_), .A3(new_n403_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT96), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n402_), .A2(new_n403_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n395_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n402_), .A2(KEYINPUT96), .A3(new_n403_), .A4(new_n395_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n419_), .A2(new_n423_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n407_), .A2(new_n421_), .A3(new_n414_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n428_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT100), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  NOR4_X1   g246(.A1(new_n431_), .A2(KEYINPUT33), .A3(new_n432_), .A4(new_n428_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n432_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n429_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n447_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n434_), .B1(new_n452_), .B2(KEYINPUT101), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT101), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n447_), .B(new_n454_), .C1(new_n451_), .C2(new_n448_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n360_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n351_), .A2(new_n359_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n433_), .A2(new_n430_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT27), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n390_), .B2(new_n439_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n435_), .A2(KEYINPUT103), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n435_), .A2(KEYINPUT103), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n442_), .A2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT104), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT104), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n442_), .A2(new_n467_), .A3(new_n460_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n459_), .A2(new_n469_), .A3(KEYINPUT105), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT105), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n442_), .A2(new_n467_), .A3(new_n460_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n442_), .B2(new_n460_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n360_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n471_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n470_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n261_), .B1(new_n456_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n469_), .A2(new_n457_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n261_), .A2(new_n458_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT106), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT106), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n469_), .A2(new_n481_), .A3(new_n484_), .A4(new_n457_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT75), .B(KEYINPUT15), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT78), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495_));
  INV_X1    g294(.A(G1gat), .ZN(new_n496_));
  INV_X1    g295(.A(G8gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT14), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n493_), .A2(KEYINPUT78), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n493_), .A2(KEYINPUT78), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n501_), .A2(new_n498_), .A3(new_n495_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n492_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n490_), .A3(new_n503_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  OR3_X1    g308(.A1(new_n505_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n490_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n504_), .A2(new_n511_), .ZN(new_n512_));
  AOI211_X1 g311(.A(KEYINPUT80), .B(new_n508_), .C1(new_n512_), .C2(new_n506_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT80), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n506_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n509_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n510_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT81), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n510_), .B(new_n523_), .C1(new_n513_), .C2(new_n516_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT82), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(KEYINPUT82), .A3(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT107), .B1(new_n487_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT107), .ZN(new_n531_));
  INV_X1    g330(.A(new_n529_), .ZN(new_n532_));
  AOI211_X1 g331(.A(new_n531_), .B(new_n532_), .C1(new_n479_), .C2(new_n486_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT74), .ZN(new_n535_));
  XOR2_X1   g334(.A(G57gat), .B(G64gat), .Z(new_n536_));
  INV_X1    g335(.A(KEYINPUT11), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT67), .B(G71gat), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G78gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT67), .B(G71gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n336_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT68), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT68), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n538_), .A2(new_n540_), .A3(new_n545_), .A4(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n536_), .A2(new_n537_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n550_), .A2(KEYINPUT71), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT71), .B1(new_n550_), .B2(new_n551_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT69), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT8), .ZN(new_n557_));
  XOR2_X1   g356(.A(G85gat), .B(G92gat), .Z(new_n558_));
  NOR2_X1   g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n557_), .B(new_n558_), .C1(new_n561_), .C2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n558_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n562_), .B(KEYINPUT6), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n561_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(KEYINPUT66), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n566_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n556_), .B(new_n565_), .C1(new_n571_), .C2(new_n557_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n567_), .ZN(new_n573_));
  OR2_X1    g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n560_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n570_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n557_), .B1(new_n576_), .B2(new_n558_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n565_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT69), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT10), .B(G99gat), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n328_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n558_), .A2(KEYINPUT9), .ZN(new_n582_));
  INV_X1    g381(.A(G85gat), .ZN(new_n583_));
  INV_X1    g382(.A(G92gat), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT9), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n581_), .A2(new_n582_), .A3(new_n585_), .A4(new_n568_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT70), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n572_), .A2(new_n579_), .A3(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n554_), .A2(new_n555_), .A3(KEYINPUT12), .A4(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n550_), .A2(new_n551_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n550_), .A2(KEYINPUT71), .A3(new_n551_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n592_), .A2(new_n588_), .A3(KEYINPUT12), .A4(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT72), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT64), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n565_), .B1(new_n571_), .B2(new_n557_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n586_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT12), .B1(new_n599_), .B2(new_n590_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n590_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n589_), .A2(new_n595_), .A3(new_n597_), .A4(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n597_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n601_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n599_), .A2(new_n590_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G120gat), .B(G148gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n603_), .A2(new_n607_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n535_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n603_), .A2(new_n607_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n612_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(KEYINPUT74), .A3(new_n614_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n620_), .A3(KEYINPUT13), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT13), .B1(new_n617_), .B2(new_n620_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n588_), .A2(new_n492_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT76), .ZN(new_n626_));
  INV_X1    g425(.A(new_n599_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT35), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT34), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n627_), .A2(new_n490_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n628_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT77), .ZN(new_n637_));
  XOR2_X1   g436(.A(G134gat), .B(G162gat), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(KEYINPUT36), .ZN(new_n641_));
  INV_X1    g440(.A(new_n634_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n626_), .A2(new_n642_), .A3(new_n632_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n635_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n639_), .B(KEYINPUT36), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n635_), .B2(new_n643_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT37), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n643_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n642_), .B1(new_n626_), .B2(new_n632_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n645_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT37), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n635_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n648_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT17), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G127gat), .B(G155gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT16), .ZN(new_n659_));
  XOR2_X1   g458(.A(G183gat), .B(G211gat), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n554_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(G231gat), .A2(G233gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n504_), .B(new_n663_), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n657_), .B(new_n661_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n664_), .B(KEYINPUT79), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(new_n590_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n590_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n661_), .B(KEYINPUT17), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n624_), .A2(new_n656_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n534_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT108), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n534_), .A2(new_n673_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT38), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n458_), .A2(new_n496_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n487_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n651_), .A2(new_n653_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n682_), .A2(new_n672_), .A3(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n624_), .A2(new_n532_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n458_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G1gat), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n679_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n681_), .A2(new_n689_), .A3(new_n690_), .ZN(G1324gat));
  OAI21_X1  g490(.A(G8gat), .B1(new_n687_), .B2(new_n469_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT39), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT39), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n694_), .B(G8gat), .C1(new_n687_), .C2(new_n469_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n475_), .A2(new_n497_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n678_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n696_), .B(KEYINPUT40), .C1(new_n678_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1325gat));
  OAI21_X1  g501(.A(G15gat), .B1(new_n687_), .B2(new_n261_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT41), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n674_), .A2(G15gat), .A3(new_n261_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1326gat));
  OAI21_X1  g505(.A(G22gat), .B1(new_n687_), .B2(new_n457_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n708_));
  XOR2_X1   g507(.A(new_n707_), .B(new_n708_), .Z(new_n709_));
  NOR3_X1   g508(.A1(new_n674_), .A2(G22gat), .A3(new_n457_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1327gat));
  NAND2_X1  g510(.A1(new_n684_), .A2(new_n672_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n624_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n713_), .B(KEYINPUT111), .C1(new_n530_), .C2(new_n533_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G29gat), .B1(new_n718_), .B2(new_n458_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n655_), .A2(KEYINPUT43), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(new_n487_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n655_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n648_), .A2(KEYINPUT110), .A3(new_n654_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n487_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n722_), .B1(new_n727_), .B2(KEYINPUT43), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n686_), .A2(new_n672_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n720_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n729_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n726_), .B2(new_n487_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n731_), .B(KEYINPUT44), .C1(new_n733_), .C2(new_n722_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n730_), .A2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n458_), .A2(G29gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n719_), .B1(new_n735_), .B2(new_n736_), .ZN(G1328gat));
  NOR2_X1   g536(.A1(new_n469_), .A2(G36gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n716_), .A2(new_n717_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT45), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n716_), .A2(new_n741_), .A3(new_n717_), .A4(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n730_), .A2(new_n734_), .A3(new_n475_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G36gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n743_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1329gat));
  INV_X1    g550(.A(new_n261_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n730_), .A2(new_n734_), .A3(G43gat), .A4(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n716_), .A2(new_n752_), .A3(new_n717_), .ZN(new_n754_));
  INV_X1    g553(.A(G43gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1330gat));
  INV_X1    g558(.A(G50gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n730_), .A2(new_n734_), .A3(new_n360_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(KEYINPUT114), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(KEYINPUT114), .B2(new_n761_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n718_), .A2(new_n760_), .A3(new_n360_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1331gat));
  OR2_X1    g564(.A1(new_n622_), .A2(new_n623_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n529_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n672_), .B1(new_n648_), .B2(new_n654_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n487_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(G57gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n458_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n685_), .A2(new_n767_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT115), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(new_n458_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n774_), .B2(new_n770_), .ZN(G1332gat));
  INV_X1    g574(.A(G64gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n776_), .A3(new_n475_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT48), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n475_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G64gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT48), .B(new_n776_), .C1(new_n773_), .C2(new_n475_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1333gat));
  NOR2_X1   g581(.A1(new_n261_), .A2(G71gat), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT116), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n769_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n773_), .A2(new_n752_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(G71gat), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT49), .B(new_n203_), .C1(new_n773_), .C2(new_n752_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1334gat));
  NAND3_X1  g589(.A1(new_n769_), .A2(new_n336_), .A3(new_n360_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n773_), .A2(new_n360_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(G78gat), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G78gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(G1335gat));
  INV_X1    g595(.A(new_n672_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n766_), .A2(new_n529_), .A3(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n733_), .B2(new_n722_), .ZN(new_n799_));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799_), .B2(new_n688_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n682_), .A2(new_n766_), .A3(new_n529_), .A4(new_n712_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n583_), .A3(new_n458_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1336gat));
  OAI21_X1  g602(.A(G92gat), .B1(new_n799_), .B2(new_n469_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n801_), .A2(new_n584_), .A3(new_n475_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n799_), .B2(new_n261_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n801_), .A2(new_n752_), .A3(new_n580_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g609(.A1(new_n801_), .A2(new_n328_), .A3(new_n360_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n798_), .B(new_n360_), .C1(new_n733_), .C2(new_n722_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(G106gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n812_), .B2(G106gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n529_), .A2(new_n614_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n603_), .A2(new_n820_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n594_), .A2(KEYINPUT72), .B1(new_n600_), .B2(new_n601_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n589_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n604_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n822_), .A2(KEYINPUT55), .A3(new_n597_), .A4(new_n589_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n612_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n819_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n505_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n509_), .B1(new_n512_), .B2(new_n506_), .ZN(new_n833_));
  OR3_X1    g632(.A1(new_n833_), .A2(KEYINPUT118), .A3(new_n523_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT118), .B1(new_n833_), .B2(new_n523_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n524_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  AOI211_X1 g637(.A(KEYINPUT119), .B(new_n832_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n617_), .A2(new_n620_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n683_), .B1(new_n831_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT57), .B(new_n683_), .C1(new_n831_), .C2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n614_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT120), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n614_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n826_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n826_), .B2(new_n612_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  OAI221_X1 g655(.A(new_n850_), .B1(new_n854_), .B2(KEYINPUT58), .C1(new_n851_), .C2(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n656_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n844_), .A2(new_n845_), .A3(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n768_), .B(new_n532_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT54), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n766_), .A2(new_n862_), .A3(new_n532_), .A4(new_n768_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n859_), .A2(new_n672_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n480_), .A2(new_n261_), .A3(new_n688_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n818_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n655_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n843_), .A2(new_n842_), .B1(new_n868_), .B2(new_n857_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n797_), .B1(new_n869_), .B2(new_n845_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n863_), .A2(new_n861_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT59), .B(new_n865_), .C1(new_n870_), .C2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n867_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n529_), .A2(G113gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT122), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n859_), .A2(new_n672_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n871_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n865_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n248_), .B1(new_n880_), .B2(new_n532_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(KEYINPUT123), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  INV_X1    g682(.A(new_n876_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n867_), .B2(new_n873_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n864_), .A2(new_n866_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G113gat), .B1(new_n886_), .B2(new_n529_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n883_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n882_), .A2(new_n888_), .ZN(G1340gat));
  OAI21_X1  g688(.A(new_n246_), .B1(new_n766_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n886_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n246_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n766_), .B1(new_n867_), .B2(new_n873_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n246_), .ZN(G1341gat));
  OAI21_X1  g692(.A(new_n243_), .B1(new_n880_), .B2(new_n672_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(KEYINPUT124), .B(new_n243_), .C1(new_n880_), .C2(new_n672_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n672_), .A2(new_n243_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n896_), .A2(new_n897_), .B1(new_n874_), .B2(new_n898_), .ZN(G1342gat));
  NAND3_X1  g698(.A1(new_n886_), .A2(new_n241_), .A3(new_n684_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n655_), .B1(new_n867_), .B2(new_n873_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n241_), .ZN(G1343gat));
  NOR4_X1   g701(.A1(new_n475_), .A2(new_n752_), .A3(new_n688_), .A4(new_n457_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n879_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n529_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT125), .B(G141gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1344gat));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n624_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n879_), .A2(new_n797_), .A3(new_n903_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT126), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n879_), .A2(new_n912_), .A3(new_n797_), .A4(new_n903_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n911_), .B2(new_n913_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1346gat));
  AOI21_X1  g716(.A(G162gat), .B1(new_n904_), .B2(new_n684_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n277_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n904_), .B2(new_n919_), .ZN(G1347gat));
  NOR3_X1   g719(.A1(new_n482_), .A2(new_n469_), .A3(new_n360_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n879_), .A2(new_n529_), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n922_), .A2(new_n923_), .A3(new_n224_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n224_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n375_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(G1348gat));
  NOR2_X1   g726(.A1(KEYINPUT127), .A2(G176gat), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n879_), .A2(new_n921_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n624_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(KEYINPUT127), .A2(G176gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  AOI211_X1 g731(.A(KEYINPUT127), .B(G176gat), .C1(new_n929_), .C2(new_n624_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1349gat));
  AOI21_X1  g733(.A(G183gat), .B1(new_n929_), .B2(new_n797_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n365_), .A2(new_n367_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n929_), .A2(new_n797_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n929_), .A2(new_n366_), .A3(new_n684_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n929_), .A2(new_n656_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n214_), .ZN(G1351gat));
  NAND3_X1  g740(.A1(new_n459_), .A2(new_n261_), .A3(new_n475_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n864_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n529_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n624_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g746(.A1(new_n864_), .A2(new_n672_), .A3(new_n942_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n948_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT63), .B(G211gat), .Z(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n948_), .B2(new_n950_), .ZN(G1354gat));
  NAND3_X1  g750(.A1(new_n943_), .A2(new_n315_), .A3(new_n684_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n864_), .A2(new_n655_), .A3(new_n942_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n315_), .ZN(G1355gat));
endmodule


