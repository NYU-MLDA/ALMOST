//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT88), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G155gat), .A3(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT1), .ZN(new_n209_));
  OR2_X1    g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n205_), .A2(new_n207_), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT87), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT89), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT2), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(KEYINPUT2), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(new_n214_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(KEYINPUT3), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n219_), .A2(new_n214_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n210_), .B(new_n208_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n217_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n217_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT91), .ZN(new_n231_));
  INV_X1    g030(.A(G204gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(G197gat), .ZN(new_n233_));
  INV_X1    g032(.A(G197gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(G197gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G211gat), .B(G218gat), .Z(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(KEYINPUT21), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(G204gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n237_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(new_n239_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(KEYINPUT21), .B2(new_n238_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT92), .A3(new_n239_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n242_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n228_), .A2(new_n230_), .A3(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n242_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n252_), .A2(new_n229_), .A3(new_n217_), .A4(new_n226_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n203_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G22gat), .B(G50gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT90), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G228gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT28), .Z(new_n259_));
  XNOR2_X1  g058(.A(new_n257_), .B(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n251_), .A2(new_n253_), .A3(new_n203_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n260_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n261_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n254_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G127gat), .ZN(new_n267_));
  INV_X1    g066(.A(G134gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G127gat), .A2(G134gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G113gat), .ZN(new_n272_));
  INV_X1    g071(.A(G113gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n273_), .A3(new_n270_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n272_), .A2(G120gat), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(G120gat), .B1(new_n272_), .B2(new_n274_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT31), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n279_));
  INV_X1    g078(.A(G169gat), .ZN(new_n280_));
  INV_X1    g079(.A(G176gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n282_), .B1(new_n285_), .B2(new_n281_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n289_));
  NAND2_X1  g088(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(KEYINPUT23), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT81), .B(G183gat), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n291_), .A2(new_n293_), .B1(G190gat), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT83), .ZN(new_n296_));
  AOI21_X1  g095(.A(G176gat), .B1(new_n283_), .B2(new_n284_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(new_n282_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G183gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT81), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G183gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n303_), .A3(KEYINPUT25), .ZN(new_n304_));
  OR2_X1    g103(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT26), .B(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n288_), .A2(KEYINPUT23), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n289_), .A2(new_n290_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n288_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n282_), .A2(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT24), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n308_), .A2(new_n313_), .A3(new_n316_), .A4(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n299_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n299_), .B2(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n279_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n299_), .A2(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT30), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n299_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n279_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G15gat), .B(G43gat), .Z(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G71gat), .B(G99gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n323_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n334_), .A2(new_n335_), .A3(KEYINPUT86), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n337_));
  INV_X1    g136(.A(new_n333_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n321_), .A2(new_n322_), .A3(new_n279_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n327_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n323_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n337_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n278_), .B1(new_n336_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n337_), .A3(new_n342_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n278_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n217_), .A2(new_n226_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n277_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n277_), .A2(new_n217_), .A3(new_n226_), .A4(new_n349_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(new_n227_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT96), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(new_n355_), .A3(new_n353_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n354_), .A2(KEYINPUT96), .A3(new_n356_), .A4(new_n358_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT0), .B(G57gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G85gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(G1gat), .B(G29gat), .Z(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT18), .B(G64gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AND4_X1   g178(.A1(KEYINPUT92), .A2(new_n238_), .A3(KEYINPUT21), .A4(new_n239_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT92), .B1(new_n248_), .B2(new_n239_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(new_n247_), .A3(new_n319_), .A4(new_n299_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT19), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n289_), .A2(new_n290_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n309_), .B1(new_n386_), .B2(new_n288_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n286_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n292_), .B1(new_n386_), .B2(new_n288_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n314_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n317_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n307_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n390_), .A2(new_n392_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n389_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n250_), .A2(new_n398_), .ZN(new_n399_));
  AND4_X1   g198(.A1(KEYINPUT20), .A2(new_n383_), .A3(new_n385_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n389_), .A2(new_n397_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n252_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n324_), .A2(new_n250_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n385_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n379_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n385_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n404_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n250_), .B2(new_n398_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n324_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n401_), .B1(new_n411_), .B2(new_n252_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n385_), .A3(new_n399_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n378_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT94), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n406_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n413_), .A2(new_n410_), .A3(KEYINPUT94), .A4(new_n378_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n368_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT33), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n354_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n352_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n368_), .A3(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n372_), .A2(new_n418_), .A3(new_n420_), .A4(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n379_), .A2(KEYINPUT32), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n385_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT97), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT97), .B(new_n385_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n383_), .A2(KEYINPUT20), .A3(new_n407_), .A4(new_n399_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT98), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n412_), .A2(KEYINPUT98), .A3(new_n407_), .A4(new_n399_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n429_), .A2(new_n430_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n362_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OAI221_X1 g236(.A(new_n426_), .B1(new_n425_), .B2(new_n435_), .C1(new_n437_), .C2(new_n419_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n348_), .B1(new_n424_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT100), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n378_), .B(KEYINPUT99), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n429_), .A2(new_n430_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n433_), .A2(new_n434_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n440_), .B(new_n442_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT100), .B1(new_n435_), .B2(new_n441_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(KEYINPUT27), .A4(new_n406_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT27), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n416_), .A2(new_n448_), .A3(new_n417_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n437_), .A2(new_n419_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n347_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT86), .B1(new_n334_), .B2(new_n335_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n346_), .B1(new_n454_), .B2(new_n345_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n266_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n262_), .A2(new_n265_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n344_), .A2(new_n457_), .A3(new_n347_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n452_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n266_), .A2(new_n439_), .B1(new_n450_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G15gat), .A2(G22gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G15gat), .A2(G22gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT76), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G15gat), .ZN(new_n466_));
  INV_X1    g265(.A(G22gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT76), .B1(new_n468_), .B2(new_n461_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G1gat), .A2(G8gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT77), .B1(new_n470_), .B2(KEYINPUT14), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n470_), .A2(KEYINPUT77), .A3(KEYINPUT14), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n465_), .A2(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G1gat), .B(G8gat), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n472_), .A2(new_n471_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n464_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n468_), .A2(KEYINPUT76), .A3(new_n461_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n474_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(G57gat), .A2(G64gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G57gat), .A2(G64gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G71gat), .B(G78gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT11), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n489_), .A3(new_n484_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n485_), .A2(new_n487_), .A3(KEYINPUT11), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n482_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT16), .B(G183gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G211gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G127gat), .B(G155gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(KEYINPUT17), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n501_), .B(KEYINPUT17), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n497_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT34), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(KEYINPUT35), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(G106gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n515_), .A2(new_n518_), .A3(new_n519_), .A4(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT8), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT8), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n521_), .A2(new_n527_), .A3(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT65), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT9), .ZN(new_n531_));
  INV_X1    g330(.A(G85gat), .ZN(new_n532_));
  INV_X1    g331(.A(G92gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n531_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n530_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n513_), .A2(KEYINPUT10), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT10), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(G99gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(G106gat), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n518_), .A2(new_n519_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(KEYINPUT65), .B(new_n537_), .C1(new_n524_), .C2(new_n531_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n511_), .B1(new_n529_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n527_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n521_), .A2(new_n527_), .A3(new_n524_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n547_), .B(new_n511_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554_));
  INV_X1    g353(.A(G43gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT72), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(G43gat), .ZN(new_n558_));
  INV_X1    g357(.A(G50gat), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G29gat), .B(G36gat), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G29gat), .B(G36gat), .Z(new_n564_));
  NOR2_X1   g363(.A1(new_n557_), .A2(G43gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n555_), .A2(KEYINPUT72), .ZN(new_n566_));
  OAI21_X1  g365(.A(G50gat), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n564_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n554_), .B1(new_n563_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n562_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(KEYINPUT15), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n510_), .B1(new_n553_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n572_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n529_), .A2(new_n577_), .A3(new_n547_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n509_), .A2(KEYINPUT35), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT71), .Z(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n552_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n575_), .B1(new_n586_), .B2(new_n548_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n510_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n587_), .A2(new_n580_), .A3(new_n588_), .A4(new_n581_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n584_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G134gat), .ZN(new_n593_));
  INV_X1    g392(.A(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT75), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n585_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n595_), .B(KEYINPUT36), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n507_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n585_), .A2(new_n591_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n600_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n585_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(KEYINPUT37), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n460_), .A2(new_n506_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT12), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n493_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n586_), .B2(new_n548_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n529_), .A2(new_n547_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n494_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n610_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n529_), .A2(new_n547_), .A3(new_n493_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT64), .Z(new_n618_));
  AND2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n615_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT66), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n616_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n529_), .A2(KEYINPUT66), .A3(new_n547_), .A4(new_n493_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(new_n614_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n620_), .B(new_n626_), .C1(new_n631_), .C2(new_n618_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n612_), .A2(new_n615_), .A3(new_n619_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n618_), .B1(new_n630_), .B2(new_n614_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n625_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n632_), .A2(new_n635_), .A3(KEYINPUT69), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT69), .B1(new_n632_), .B2(new_n635_), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n636_), .A2(new_n637_), .B1(KEYINPUT70), .B2(KEYINPUT13), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n635_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT69), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n635_), .A3(KEYINPUT69), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n638_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n474_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n473_), .A2(new_n475_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n570_), .B(new_n573_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G229gat), .A2(G233gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n476_), .A2(new_n577_), .A3(new_n481_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n650_), .A2(KEYINPUT78), .A3(new_n651_), .A4(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(new_n280_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(G197gat), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT78), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n572_), .B(new_n571_), .C1(new_n649_), .C2(new_n648_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n652_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n651_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n653_), .B(new_n656_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT79), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n651_), .B1(new_n658_), .B2(new_n652_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n650_), .A2(new_n652_), .ZN(new_n666_));
  OAI22_X1  g465(.A1(new_n665_), .A2(new_n657_), .B1(new_n666_), .B2(new_n660_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n656_), .B1(new_n667_), .B2(new_n653_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT79), .B(new_n656_), .C1(new_n667_), .C2(new_n653_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(KEYINPUT80), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT80), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n664_), .A2(new_n668_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n670_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n647_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n609_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(G1gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n452_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT38), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n599_), .A2(new_n602_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n460_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n674_), .A2(new_n670_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n506_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n646_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT101), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT101), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G1gat), .B1(new_n689_), .B2(new_n451_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n681_), .A2(new_n690_), .ZN(G1324gat));
  INV_X1    g490(.A(G8gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n450_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n678_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G8gat), .B1(new_n689_), .B2(new_n450_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT39), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT40), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n696_), .A2(KEYINPUT40), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1325gat));
  INV_X1    g502(.A(new_n348_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G15gat), .B1(new_n689_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT104), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n705_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n678_), .A2(new_n466_), .A3(new_n348_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT105), .ZN(G1326gat));
  OAI21_X1  g510(.A(G22gat), .B1(new_n689_), .B2(new_n266_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT42), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n678_), .A2(new_n467_), .A3(new_n457_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1327gat));
  NAND2_X1  g514(.A1(new_n424_), .A2(new_n438_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n266_), .A3(new_n704_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n456_), .A2(new_n458_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n718_), .A2(new_n451_), .A3(new_n449_), .A4(new_n447_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n720_), .A2(new_n682_), .A3(new_n677_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(new_n506_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G29gat), .B1(new_n722_), .B2(new_n452_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n603_), .A2(new_n607_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n726_), .A3(new_n608_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n646_), .A2(new_n684_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n506_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n728_), .A2(KEYINPUT44), .A3(new_n729_), .A4(new_n506_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n452_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n723_), .B1(new_n734_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n693_), .A3(new_n733_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G36gat), .ZN(new_n737_));
  INV_X1    g536(.A(G36gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n722_), .A2(new_n738_), .A3(new_n693_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT45), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n740_), .A3(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  NAND3_X1  g544(.A1(new_n732_), .A2(new_n348_), .A3(new_n733_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G43gat), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n722_), .A2(new_n555_), .A3(new_n348_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1330gat));
  NAND3_X1  g551(.A1(new_n732_), .A2(new_n457_), .A3(new_n733_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n754_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(G50gat), .A3(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n722_), .A2(new_n559_), .A3(new_n457_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1331gat));
  NOR2_X1   g558(.A1(new_n646_), .A2(new_n684_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n609_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n452_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n506_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n683_), .A2(new_n647_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(new_n451_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n762_), .B1(new_n766_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g566(.A(G64gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n764_), .B2(new_n693_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT48), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n761_), .A2(new_n768_), .A3(new_n693_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1333gat));
  NOR2_X1   g571(.A1(new_n704_), .A2(G71gat), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT107), .Z(new_n774_));
  NAND2_X1  g573(.A1(new_n761_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n764_), .A2(new_n348_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G71gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G71gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1334gat));
  OAI21_X1  g581(.A(G78gat), .B1(new_n765_), .B2(new_n266_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n783_), .A2(KEYINPUT109), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT109), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(G78gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n761_), .A2(new_n789_), .A3(new_n457_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n784_), .A2(KEYINPUT50), .A3(new_n785_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(new_n790_), .A3(new_n791_), .ZN(G1335gat));
  NOR3_X1   g591(.A1(new_n646_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n720_), .A2(new_n682_), .A3(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT110), .Z(new_n795_));
  AOI21_X1  g594(.A(G85gat), .B1(new_n795_), .B2(new_n452_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT111), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n728_), .A2(new_n793_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(G85gat), .A3(new_n452_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1336gat));
  AOI21_X1  g599(.A(G92gat), .B1(new_n795_), .B2(new_n693_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n450_), .A2(new_n533_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT112), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n798_), .B2(new_n803_), .ZN(G1337gat));
  NAND2_X1  g603(.A1(new_n540_), .A2(new_n542_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n795_), .A2(new_n805_), .A3(new_n348_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n513_), .B1(new_n798_), .B2(new_n348_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g608(.A(new_n726_), .B1(new_n720_), .B2(new_n608_), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT43), .B(new_n724_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n457_), .B(new_n793_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT113), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n728_), .A2(new_n814_), .A3(new_n457_), .A4(new_n793_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n815_), .A3(G106gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n813_), .A2(new_n815_), .A3(G106gat), .A4(new_n817_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n795_), .A2(new_n514_), .A3(new_n457_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT53), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n825_), .A3(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1339gat));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n608_), .B1(new_n645_), .B2(new_n638_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n763_), .ZN(new_n830_));
  AND4_X1   g629(.A1(new_n828_), .A2(new_n763_), .A3(new_n646_), .A4(new_n724_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n666_), .A2(KEYINPUT115), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n666_), .A2(KEYINPUT115), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n660_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n656_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n659_), .A2(new_n651_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n663_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n612_), .A2(new_n630_), .A3(new_n615_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n618_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n620_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n612_), .A2(new_n615_), .A3(KEYINPUT55), .A4(new_n619_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n625_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n848_), .B2(new_n625_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n632_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n841_), .B1(new_n853_), .B2(new_n684_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT116), .B(new_n833_), .C1(new_n854_), .C2(new_n682_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n625_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT56), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n848_), .A2(new_n849_), .A3(new_n625_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n684_), .A2(new_n857_), .A3(new_n632_), .A4(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n840_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n682_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT57), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n853_), .A2(KEYINPUT58), .A3(new_n860_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n857_), .A2(new_n632_), .A3(new_n858_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n840_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n868_), .A3(new_n608_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n855_), .A2(new_n864_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n832_), .B1(new_n870_), .B2(new_n506_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n693_), .A2(new_n451_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n871_), .A2(new_n456_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G113gat), .B1(new_n874_), .B2(new_n684_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n506_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n832_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n456_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT59), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n871_), .A2(new_n881_), .A3(new_n456_), .A4(new_n873_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n273_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n676_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n875_), .B1(new_n884_), .B2(new_n885_), .ZN(G1340gat));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT117), .B(G120gat), .Z(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n876_), .A2(new_n877_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n879_), .A3(new_n872_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n881_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n878_), .A2(KEYINPUT59), .A3(new_n879_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n889_), .B1(new_n894_), .B2(new_n647_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n889_), .B1(new_n646_), .B2(KEYINPUT60), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n889_), .A2(KEYINPUT60), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n878_), .A2(new_n879_), .A3(new_n896_), .A4(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n874_), .A2(KEYINPUT118), .A3(new_n896_), .A4(new_n897_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n887_), .B1(new_n895_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n888_), .B1(new_n883_), .B2(new_n646_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n901_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(KEYINPUT119), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(G1341gat));
  OAI21_X1  g706(.A(new_n267_), .B1(new_n891_), .B2(new_n506_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT120), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n883_), .A2(new_n506_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(G127gat), .B2(new_n910_), .ZN(G1342gat));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n608_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G134gat), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n682_), .A2(new_n268_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n891_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n912_), .B1(new_n914_), .B2(new_n917_), .ZN(new_n918_));
  AOI211_X1 g717(.A(KEYINPUT121), .B(new_n916_), .C1(new_n913_), .C2(G134gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1343gat));
  NOR3_X1   g719(.A1(new_n871_), .A2(new_n458_), .A3(new_n873_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n684_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n647_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n685_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT61), .B(G155gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n921_), .B2(new_n682_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n921_), .A2(new_n608_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(G162gat), .B2(new_n930_), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n871_), .A2(new_n456_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n450_), .A2(new_n452_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n684_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(G169gat), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n940_));
  INV_X1    g739(.A(new_n285_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n939_), .B(new_n940_), .C1(new_n941_), .C2(new_n936_), .ZN(G1348gat));
  XOR2_X1   g741(.A(KEYINPUT122), .B(G176gat), .Z(new_n943_));
  NAND3_X1  g742(.A1(new_n935_), .A2(new_n647_), .A3(new_n943_), .ZN(new_n944_));
  OAI22_X1  g743(.A1(new_n934_), .A2(new_n646_), .B1(KEYINPUT122), .B2(new_n281_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1349gat));
  NAND2_X1  g745(.A1(new_n935_), .A2(new_n685_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n294_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n395_), .B1(new_n294_), .B2(KEYINPUT123), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n947_), .B2(new_n950_), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n935_), .A2(new_n682_), .A3(new_n307_), .ZN(new_n952_));
  OAI21_X1  g751(.A(G190gat), .B1(new_n934_), .B2(new_n724_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1351gat));
  NOR2_X1   g753(.A1(new_n871_), .A2(new_n458_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n933_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n957_), .A2(G197gat), .A3(new_n684_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n958_), .A2(KEYINPUT124), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(KEYINPUT124), .ZN(new_n960_));
  AOI21_X1  g759(.A(G197gat), .B1(new_n957_), .B2(new_n684_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(G1352gat));
  OR2_X1    g761(.A1(new_n232_), .A2(KEYINPUT125), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n957_), .A2(new_n647_), .A3(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n232_), .A2(KEYINPUT125), .ZN(new_n965_));
  XOR2_X1   g764(.A(new_n965_), .B(KEYINPUT126), .Z(new_n966_));
  XOR2_X1   g765(.A(new_n964_), .B(new_n966_), .Z(G1353gat));
  NOR2_X1   g766(.A1(new_n956_), .A2(new_n506_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n968_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969_));
  XOR2_X1   g768(.A(KEYINPUT63), .B(G211gat), .Z(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(new_n968_), .B2(new_n970_), .ZN(G1354gat));
  INV_X1    g770(.A(new_n682_), .ZN(new_n972_));
  OR3_X1    g771(.A1(new_n956_), .A2(KEYINPUT127), .A3(new_n972_), .ZN(new_n973_));
  INV_X1    g772(.A(G218gat), .ZN(new_n974_));
  OAI21_X1  g773(.A(KEYINPUT127), .B1(new_n956_), .B2(new_n972_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n973_), .A2(new_n974_), .A3(new_n975_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n957_), .A2(G218gat), .A3(new_n608_), .ZN(new_n977_));
  AND2_X1   g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1355gat));
endmodule


