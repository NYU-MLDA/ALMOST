//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_;
  INV_X1    g000(.A(G190gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT26), .B1(new_n202_), .B2(KEYINPUT82), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT82), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT26), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G183gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n213_), .A2(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT83), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT83), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G169gat), .A3(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n211_), .A2(new_n218_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n222_), .A2(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n212_), .A2(new_n214_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n207_), .A2(new_n202_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT22), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n228_), .A2(new_n232_), .A3(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n226_), .A2(new_n227_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n227_), .B1(new_n226_), .B2(new_n239_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G99gat), .ZN(new_n243_));
  INV_X1    g042(.A(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n242_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT85), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT85), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n247_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n246_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(G15gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT30), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT31), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G8gat), .B(G36gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G197gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G204gat), .ZN(new_n272_));
  INV_X1    g071(.A(G204gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G197gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT21), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n273_), .B2(G197gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .A4(new_n274_), .ZN(new_n281_));
  INV_X1    g080(.A(G218gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G211gat), .ZN(new_n283_));
  INV_X1    g082(.A(G211gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G218gat), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n276_), .A2(new_n281_), .A3(new_n283_), .A4(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n278_), .A2(new_n279_), .A3(new_n274_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n280_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n289_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n286_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n240_), .A2(new_n292_), .A3(new_n241_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT20), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT90), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT19), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n287_), .A2(new_n288_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT88), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n283_), .A2(new_n285_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(KEYINPUT21), .B2(new_n275_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n300_), .A2(new_n301_), .B1(new_n281_), .B2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n228_), .A2(new_n238_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n208_), .A2(new_n210_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT26), .B(G190gat), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n306_), .A2(new_n307_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n305_), .A2(new_n232_), .B1(new_n308_), .B2(new_n218_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n226_), .A2(new_n239_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT84), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n226_), .A2(new_n227_), .A3(new_n239_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n304_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(KEYINPUT20), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n295_), .A2(new_n298_), .A3(new_n311_), .A4(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT97), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n308_), .A2(new_n218_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n239_), .ZN(new_n322_));
  OAI211_X1 g121(.A(KEYINPUT96), .B(new_n320_), .C1(new_n322_), .C2(new_n292_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n292_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n304_), .A2(new_n309_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT96), .B1(new_n326_), .B2(new_n320_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n319_), .B(new_n297_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n318_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n320_), .B1(new_n322_), .B2(new_n292_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT96), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n324_), .A3(new_n323_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n319_), .B1(new_n333_), .B2(new_n297_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n270_), .B1(new_n329_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT98), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n317_), .A2(new_n311_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n316_), .B1(new_n315_), .B2(KEYINPUT20), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n297_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n324_), .A2(KEYINPUT20), .A3(new_n298_), .A4(new_n326_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n270_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT99), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n340_), .A2(KEYINPUT99), .A3(new_n270_), .A4(new_n341_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n336_), .A2(new_n337_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT27), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n318_), .A2(new_n328_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n269_), .B1(new_n348_), .B2(new_n334_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n349_), .B2(KEYINPUT98), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n342_), .A2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n340_), .A2(KEYINPUT92), .A3(new_n270_), .A4(new_n341_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n340_), .A2(new_n341_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n269_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n346_), .A2(new_n350_), .B1(new_n347_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G233gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n358_), .A2(KEYINPUT86), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(KEYINPUT86), .ZN(new_n360_));
  OAI21_X1  g159(.A(G228gat), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n365_), .B(KEYINPUT3), .Z(new_n366_));
  NAND2_X1  g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT2), .Z(new_n368_));
  OAI211_X1 g167(.A(new_n362_), .B(new_n364_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n363_), .B1(KEYINPUT1), .B2(new_n362_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(KEYINPUT1), .B2(new_n362_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n365_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n361_), .B1(new_n376_), .B2(new_n292_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(KEYINPUT29), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n378_), .A2(new_n361_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n292_), .B2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G78gat), .B(G106gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n374_), .A2(KEYINPUT29), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT28), .ZN(new_n384_));
  XOR2_X1   g183(.A(G22gat), .B(G50gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n382_), .B(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n255_), .A2(new_n374_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n250_), .A2(new_n254_), .A3(new_n369_), .A4(new_n373_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G1gat), .B(G29gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT93), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n390_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n255_), .A2(new_n374_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n393_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n395_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n401_), .B1(new_n395_), .B2(new_n405_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n387_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n357_), .A2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n348_), .B2(new_n334_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(KEYINPUT94), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n408_), .B(new_n412_), .C1(new_n354_), .C2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n392_), .A2(new_n394_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n402_), .A2(new_n393_), .A3(new_n404_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n400_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT33), .ZN(new_n418_));
  MUX2_X1   g217(.A(KEYINPUT33), .B(new_n418_), .S(new_n407_), .Z(new_n419_));
  OAI21_X1  g218(.A(new_n414_), .B1(new_n419_), .B2(new_n356_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n387_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n264_), .B1(new_n410_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n408_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n264_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n344_), .A2(new_n345_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n349_), .A2(KEYINPUT98), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n337_), .B(new_n269_), .C1(new_n348_), .C2(new_n334_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT27), .A4(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n356_), .A2(new_n347_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n387_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT100), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT100), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n428_), .A2(new_n429_), .A3(new_n387_), .A4(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n424_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n422_), .B1(new_n423_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n436_), .B(KEYINPUT6), .Z(new_n437_));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n440_), .A2(new_n441_), .B1(G99gat), .B2(G106gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT68), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n437_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n446_), .B2(new_n445_), .ZN(new_n448_));
  INV_X1    g247(.A(G85gat), .ZN(new_n449_));
  INV_X1    g248(.A(G92gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G85gat), .A2(G92gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n448_), .A2(KEYINPUT8), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT8), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n445_), .B2(new_n437_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n451_), .B2(KEYINPUT9), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n451_), .A2(KEYINPUT9), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n451_), .A2(KEYINPUT66), .A3(KEYINPUT9), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT10), .B(G99gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT65), .B(G106gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n437_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n455_), .A2(new_n456_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n454_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT70), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G29gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT71), .ZN(new_n471_));
  XOR2_X1   g270(.A(G43gat), .B(G50gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n454_), .A2(KEYINPUT70), .A3(new_n466_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n469_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n467_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n473_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G232gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT34), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n481_), .A2(KEYINPUT35), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(KEYINPUT35), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n477_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT75), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT75), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n477_), .A2(new_n487_), .A3(new_n479_), .A4(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n477_), .A2(new_n479_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT73), .B1(new_n490_), .B2(new_n482_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n490_), .A2(KEYINPUT73), .A3(new_n482_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT76), .ZN(new_n494_));
  XOR2_X1   g293(.A(G190gat), .B(G218gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(G134gat), .B(G162gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n493_), .B2(KEYINPUT76), .ZN(new_n500_));
  INV_X1    g299(.A(new_n491_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n490_), .A2(KEYINPUT73), .A3(new_n482_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n501_), .A2(new_n502_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n498_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT74), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n494_), .A2(new_n500_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT77), .B(G15gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G22gat), .ZN(new_n508_));
  INV_X1    g307(.A(G1gat), .ZN(new_n509_));
  INV_X1    g308(.A(G8gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT14), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G1gat), .B(G8gat), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n513_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT78), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G231gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT11), .Z(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT69), .B(G71gat), .ZN(new_n522_));
  INV_X1    g321(.A(G78gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n519_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G127gat), .B(G155gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT16), .ZN(new_n532_));
  XOR2_X1   g331(.A(G183gat), .B(G211gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n534_), .B(KEYINPUT80), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT17), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n530_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n435_), .A2(new_n506_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n478_), .A2(new_n529_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n467_), .A2(new_n528_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G230gat), .A2(G233gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT64), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n469_), .A2(KEYINPUT12), .A3(new_n528_), .A4(new_n476_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n478_), .B2(new_n529_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n544_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G120gat), .B(G148gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G176gat), .B(G204gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n554_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT13), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n516_), .B(new_n473_), .Z(new_n562_));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n475_), .A2(new_n516_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n514_), .A2(new_n473_), .A3(new_n515_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n566_), .A2(new_n563_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n562_), .A2(new_n564_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT81), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G169gat), .B(G197gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n568_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n561_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n542_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(G1gat), .B1(new_n576_), .B2(new_n423_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT103), .Z(new_n578_));
  NOR2_X1   g377(.A1(new_n435_), .A2(new_n574_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n537_), .A2(new_n540_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n503_), .A2(new_n499_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n503_), .A2(new_n505_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT37), .A3(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n580_), .B(new_n583_), .C1(new_n506_), .C2(KEYINPUT37), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n561_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n408_), .B(KEYINPUT101), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n586_), .A2(G1gat), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n578_), .A2(new_n591_), .ZN(G1324gat));
  INV_X1    g391(.A(new_n357_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n579_), .A2(new_n510_), .A3(new_n593_), .A4(new_n585_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  INV_X1    g394(.A(new_n576_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n593_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n597_), .B2(G8gat), .ZN(new_n598_));
  AOI211_X1 g397(.A(KEYINPUT39), .B(new_n510_), .C1(new_n596_), .C2(new_n593_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n594_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(G1325gat));
  OAI21_X1  g401(.A(G15gat), .B1(new_n576_), .B2(new_n424_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(KEYINPUT104), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT104), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n604_), .A2(KEYINPUT41), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT41), .B1(new_n604_), .B2(new_n605_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n586_), .A2(G15gat), .A3(new_n424_), .ZN(new_n608_));
  OR3_X1    g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(G1326gat));
  OAI21_X1  g408(.A(G22gat), .B1(new_n576_), .B2(new_n387_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT42), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n387_), .A2(G22gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n586_), .B2(new_n612_), .ZN(G1327gat));
  INV_X1    g412(.A(KEYINPUT106), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n506_), .A2(new_n541_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n561_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n579_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n431_), .A2(new_n433_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n423_), .A3(new_n264_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n422_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n573_), .A3(new_n616_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT106), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n617_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(G29gat), .B1(new_n624_), .B2(new_n408_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT43), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n583_), .B1(new_n506_), .B2(KEYINPUT37), .ZN(new_n627_));
  AOI211_X1 g426(.A(new_n408_), .B(new_n424_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n626_), .B(new_n627_), .C1(new_n628_), .C2(new_n422_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT105), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n621_), .A2(new_n631_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n627_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT43), .B1(new_n435_), .B2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n630_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n561_), .A2(new_n580_), .A3(new_n574_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n635_), .A2(KEYINPUT44), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT44), .B1(new_n635_), .B2(new_n636_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n587_), .A2(G29gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n625_), .B1(new_n639_), .B2(new_n640_), .ZN(G1328gat));
  INV_X1    g440(.A(G36gat), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n357_), .A2(KEYINPUT107), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n357_), .A2(KEYINPUT107), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n617_), .A2(new_n623_), .A3(new_n642_), .A4(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT45), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n637_), .A2(new_n638_), .A3(new_n357_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(new_n642_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n647_), .B(KEYINPUT46), .C1(new_n648_), .C2(new_n642_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1329gat));
  NAND3_X1  g452(.A1(new_n617_), .A2(new_n623_), .A3(new_n264_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n244_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NOR4_X1   g456(.A1(new_n637_), .A2(new_n638_), .A3(new_n244_), .A4(new_n424_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT47), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n639_), .A2(G43gat), .A3(new_n264_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n655_), .B(KEYINPUT108), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n663_), .ZN(G1330gat));
  INV_X1    g463(.A(new_n387_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G50gat), .B1(new_n624_), .B2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(G50gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n639_), .B2(new_n667_), .ZN(G1331gat));
  NOR2_X1   g467(.A1(new_n560_), .A2(new_n573_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n542_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(G57gat), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n423_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT109), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n435_), .A2(new_n573_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n584_), .A2(new_n560_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n671_), .B1(new_n677_), .B2(new_n588_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(KEYINPUT109), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n674_), .A2(new_n678_), .A3(new_n679_), .ZN(G1332gat));
  INV_X1    g479(.A(new_n645_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G64gat), .B1(new_n670_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT48), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n681_), .A2(G64gat), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT110), .Z(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n677_), .B2(new_n685_), .ZN(G1333gat));
  OAI21_X1  g485(.A(G71gat), .B1(new_n670_), .B2(new_n424_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n424_), .A2(G71gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n677_), .B2(new_n690_), .ZN(G1334gat));
  OAI21_X1  g490(.A(G78gat), .B1(new_n670_), .B2(new_n387_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT50), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n387_), .A2(G78gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT112), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n677_), .B2(new_n695_), .ZN(G1335gat));
  NAND4_X1  g495(.A1(new_n675_), .A2(new_n561_), .A3(new_n506_), .A4(new_n541_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT113), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n449_), .B1(new_n699_), .B2(new_n588_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n669_), .A2(new_n541_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT114), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n408_), .A2(G85gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT115), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n635_), .A2(new_n702_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT116), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n700_), .A2(KEYINPUT116), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1336gat));
  NAND2_X1  g509(.A1(new_n635_), .A2(new_n702_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G92gat), .B1(new_n711_), .B2(new_n681_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n593_), .A2(new_n450_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n699_), .B2(new_n713_), .ZN(G1337gat));
  OAI21_X1  g513(.A(G99gat), .B1(new_n711_), .B2(new_n424_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n264_), .A2(new_n463_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n699_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g517(.A(new_n697_), .B(KEYINPUT113), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n464_), .A3(new_n665_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n635_), .A2(new_n665_), .A3(new_n702_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(G106gat), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G106gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT53), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n720_), .B(new_n727_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1339gat));
  AOI21_X1  g528(.A(new_n572_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n565_), .A2(new_n566_), .A3(new_n564_), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n568_), .A2(new_n572_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n559_), .A2(new_n732_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n554_), .A2(new_n558_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n553_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n549_), .A2(new_n543_), .A3(new_n552_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n547_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT55), .A4(new_n552_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n740_), .B2(new_n558_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n573_), .B(new_n734_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n506_), .B1(new_n733_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT119), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n741_), .A2(new_n742_), .A3(KEYINPUT118), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n740_), .A2(new_n558_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(KEYINPUT118), .A3(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n734_), .A2(new_n732_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n747_), .B1(new_n748_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  INV_X1    g554(.A(new_n742_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n734_), .A2(new_n732_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n742_), .B2(KEYINPUT118), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n761_), .A3(KEYINPUT119), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n754_), .A2(new_n755_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT120), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n627_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(new_n761_), .A3(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n763_), .B2(new_n627_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n746_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n541_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n585_), .B2(new_n574_), .ZN(new_n772_));
  NOR4_X1   g571(.A1(new_n584_), .A2(KEYINPUT54), .A3(new_n573_), .A4(new_n561_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n434_), .A2(new_n587_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(KEYINPUT59), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n774_), .B1(new_n769_), .B2(new_n541_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n777_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n573_), .A2(G113gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT121), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n573_), .A3(new_n778_), .ZN(new_n786_));
  INV_X1    g585(.A(G113gat), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n783_), .A2(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(G1340gat));
  AOI21_X1  g587(.A(new_n560_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n789_));
  INV_X1    g588(.A(G120gat), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n776_), .A2(new_n778_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n560_), .B2(KEYINPUT60), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(KEYINPUT60), .B2(new_n790_), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n789_), .A2(new_n790_), .B1(new_n791_), .B2(new_n793_), .ZN(G1341gat));
  INV_X1    g593(.A(G127gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n580_), .B2(KEYINPUT122), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(KEYINPUT122), .B2(new_n795_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n776_), .A2(new_n580_), .A3(new_n778_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n783_), .A2(new_n797_), .B1(new_n798_), .B2(new_n795_), .ZN(G1342gat));
  INV_X1    g598(.A(G134gat), .ZN(new_n800_));
  INV_X1    g599(.A(new_n506_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT123), .B(new_n800_), .C1(new_n791_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT123), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n781_), .A2(new_n801_), .A3(new_n777_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(G134gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n627_), .A2(G134gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT124), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n802_), .A2(new_n805_), .B1(new_n783_), .B2(new_n807_), .ZN(G1343gat));
  NAND4_X1  g607(.A1(new_n681_), .A2(new_n665_), .A3(new_n424_), .A4(new_n587_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT125), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n776_), .A2(new_n573_), .A3(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g611(.A1(new_n776_), .A2(new_n561_), .A3(new_n810_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g613(.A1(new_n776_), .A2(new_n580_), .A3(new_n810_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1346gat));
  AND2_X1   g616(.A1(new_n776_), .A2(new_n810_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n506_), .ZN(new_n819_));
  INV_X1    g618(.A(G162gat), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n627_), .A2(G162gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT126), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n819_), .A2(new_n820_), .B1(new_n818_), .B2(new_n822_), .ZN(G1347gat));
  NOR4_X1   g622(.A1(new_n681_), .A2(new_n665_), .A3(new_n424_), .A4(new_n587_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n781_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT62), .B(G169gat), .C1(new_n827_), .C2(new_n574_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n781_), .A2(new_n574_), .A3(new_n825_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n233_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n831_), .A3(new_n832_), .ZN(G1348gat));
  NAND2_X1  g632(.A1(new_n826_), .A2(new_n561_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g634(.A1(new_n827_), .A2(new_n306_), .A3(new_n541_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G183gat), .B1(new_n826_), .B2(new_n580_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1350gat));
  OAI21_X1  g637(.A(G190gat), .B1(new_n827_), .B2(new_n633_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n307_), .A3(new_n506_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1351gat));
  NAND3_X1  g640(.A1(new_n645_), .A2(new_n409_), .A3(new_n424_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n770_), .B2(new_n775_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n573_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n561_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g646(.A1(new_n781_), .A2(new_n541_), .A3(new_n842_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT63), .B(G211gat), .Z(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n848_), .B2(new_n850_), .ZN(G1354gat));
  AOI21_X1  g650(.A(new_n282_), .B1(new_n843_), .B2(new_n627_), .ZN(new_n852_));
  NOR4_X1   g651(.A1(new_n781_), .A2(G218gat), .A3(new_n801_), .A4(new_n842_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT127), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n843_), .A2(new_n282_), .A3(new_n506_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT127), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n781_), .A2(new_n633_), .A3(new_n842_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n855_), .B(new_n856_), .C1(new_n857_), .C2(new_n282_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(G1355gat));
endmodule


