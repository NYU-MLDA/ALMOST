//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_;
  XNOR2_X1  g000(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT102), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT25), .B(G183gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT23), .Z(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n209_), .B1(new_n210_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n220_), .A2(KEYINPUT83), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(KEYINPUT83), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n207_), .B(new_n217_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n209_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT84), .B(G176gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G169gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n218_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n230_), .B(new_n233_), .Z(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G134gat), .Z(new_n235_));
  XOR2_X1   g034(.A(G113gat), .B(G120gat), .Z(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  XOR2_X1   g036(.A(new_n234_), .B(new_n237_), .Z(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n238_), .B(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G8gat), .B(G36gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G64gat), .B(G92gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT19), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT20), .ZN(new_n254_));
  XOR2_X1   g053(.A(G197gat), .B(G204gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT87), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(G204gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT21), .B(new_n262_), .C1(new_n255_), .C2(new_n260_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n263_), .B(new_n257_), .C1(KEYINPUT21), .C2(new_n255_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n254_), .B1(new_n230_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n228_), .A2(new_n218_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n267_), .A2(KEYINPUT90), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(KEYINPUT90), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n225_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT91), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n216_), .B1(new_n273_), .B2(new_n219_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(new_n273_), .B2(new_n219_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n207_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT89), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(KEYINPUT89), .A3(new_n207_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n217_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n270_), .A2(new_n271_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n253_), .B(new_n266_), .C1(new_n282_), .C2(new_n265_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT92), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n230_), .B2(new_n265_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n282_), .B2(new_n265_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n286_), .B2(new_n253_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(new_n284_), .A3(new_n253_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n250_), .B(new_n283_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n266_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n265_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n280_), .A2(new_n292_), .A3(new_n270_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n252_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT96), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n294_), .A2(new_n295_), .B1(new_n286_), .B2(new_n253_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT96), .B(new_n252_), .C1(new_n291_), .C2(new_n293_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n250_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT97), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n290_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n295_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n286_), .A2(new_n253_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n249_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT27), .B1(new_n304_), .B2(KEYINPUT97), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT98), .B1(new_n300_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT98), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(KEYINPUT97), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .A4(new_n290_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n285_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n272_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n292_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(KEYINPUT92), .A3(new_n252_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n287_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n250_), .B1(new_n317_), .B2(new_n283_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n283_), .ZN(new_n319_));
  AOI211_X1 g118(.A(new_n249_), .B(new_n319_), .C1(new_n316_), .C2(new_n287_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n307_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT99), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT99), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n323_), .B(new_n307_), .C1(new_n318_), .C2(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G155gat), .ZN(new_n326_));
  INV_X1    g125(.A(G162gat), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT1), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT1), .B1(new_n326_), .B2(new_n327_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n328_), .B(new_n329_), .C1(G155gat), .C2(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  OR2_X1    g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT85), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(KEYINPUT3), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n332_), .A2(KEYINPUT3), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n331_), .A2(new_n340_), .ZN(new_n341_));
  NOR4_X1   g140(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .A4(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n333_), .B1(new_n335_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(KEYINPUT29), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT28), .Z(new_n345_));
  AOI21_X1  g144(.A(new_n292_), .B1(KEYINPUT29), .B2(new_n343_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(G78gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G106gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G22gat), .B(G50gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n347_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  OR2_X1    g158(.A1(new_n343_), .A2(new_n237_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n343_), .A2(new_n237_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(KEYINPUT4), .A3(new_n361_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n361_), .A2(KEYINPUT4), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n359_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n365_), .A2(new_n368_), .A3(new_n359_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n355_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n312_), .A2(new_n325_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n317_), .A2(new_n283_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n249_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n369_), .A2(KEYINPUT33), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n369_), .A2(KEYINPUT33), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n359_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n366_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT94), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(KEYINPUT94), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n378_), .A2(new_n379_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n377_), .A2(new_n385_), .A3(new_n290_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT95), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n250_), .A2(KEYINPUT32), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n372_), .B1(new_n303_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n376_), .B2(new_n389_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n377_), .A2(new_n385_), .A3(KEYINPUT95), .A4(new_n290_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n355_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n244_), .B1(new_n375_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n312_), .A2(new_n325_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n355_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n244_), .A2(new_n372_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G29gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT71), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G43gat), .B(G50gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n401_), .A2(KEYINPUT71), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(KEYINPUT71), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G15gat), .B(G22gat), .ZN(new_n410_));
  INV_X1    g209(.A(G1gat), .ZN(new_n411_));
  INV_X1    g210(.A(G8gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT14), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G8gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n409_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G229gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n409_), .B(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(new_n416_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n409_), .A2(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n418_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n420_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G113gat), .B(G141gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT80), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G169gat), .B(G197gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n428_), .B(new_n429_), .Z(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n430_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n420_), .B(new_n432_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT81), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n400_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n437_));
  INV_X1    g236(.A(G99gat), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(new_n351_), .A3(KEYINPUT66), .A4(KEYINPUT7), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT64), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT64), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT6), .ZN(new_n447_));
  AND2_X1   g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n446_), .A2(KEYINPUT6), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n444_), .A2(KEYINPUT64), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n443_), .A2(new_n449_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G85gat), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n457_), .A2(KEYINPUT67), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n437_), .B1(new_n454_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n454_), .A2(new_n437_), .A3(new_n459_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n453_), .A2(new_n449_), .ZN(new_n464_));
  OR2_X1    g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n351_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(KEYINPUT9), .A3(new_n458_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n458_), .A2(KEYINPUT9), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n463_), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n445_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n448_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n472_), .A2(new_n475_), .A3(KEYINPUT65), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n461_), .A2(new_n462_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G57gat), .B(G64gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n477_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n477_), .A2(new_n484_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(G230gat), .A2(G233gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n488_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n454_), .A2(new_n437_), .A3(new_n459_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n464_), .A2(new_n470_), .A3(new_n463_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT65), .B1(new_n472_), .B2(new_n475_), .ZN(new_n495_));
  OAI22_X1  g294(.A1(new_n493_), .A2(new_n460_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT69), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n476_), .A2(new_n471_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT69), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n498_), .B(new_n499_), .C1(new_n460_), .C2(new_n493_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n481_), .B(KEYINPUT12), .C1(new_n482_), .C2(new_n483_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n477_), .B2(new_n484_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n490_), .B1(new_n477_), .B2(new_n484_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n492_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G120gat), .B(G148gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT5), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G176gat), .B(G204gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n492_), .A2(new_n507_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(KEYINPUT13), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n436_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n422_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT73), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT73), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n422_), .A2(new_n497_), .A3(new_n525_), .A4(new_n500_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n477_), .A2(new_n408_), .A3(new_n405_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT34), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT35), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n527_), .B2(KEYINPUT74), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(KEYINPUT35), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n527_), .B(new_n528_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n528_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n527_), .A2(KEYINPUT74), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n531_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G190gat), .B(G218gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n543_), .B(KEYINPUT36), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n545_), .B(KEYINPUT37), .C1(new_n538_), .C2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT77), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n538_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n534_), .A2(new_n537_), .A3(KEYINPUT77), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n550_), .A2(new_n551_), .B1(new_n544_), .B2(new_n538_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n548_), .B1(new_n552_), .B2(KEYINPUT37), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n484_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT78), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n416_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558_));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(KEYINPUT17), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n553_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT79), .ZN(new_n569_));
  NOR4_X1   g368(.A1(new_n522_), .A2(G1gat), .A3(new_n372_), .A4(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n202_), .A2(new_n203_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n204_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT101), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n306_), .A2(new_n311_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n574_), .A2(new_n374_), .B1(new_n393_), .B2(new_n355_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n355_), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n575_), .A2(new_n244_), .B1(new_n576_), .B2(new_n398_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n552_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n573_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n573_), .B(new_n578_), .C1(new_n395_), .C2(new_n399_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n434_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n567_), .A2(new_n520_), .A3(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n582_), .A2(new_n373_), .A3(new_n584_), .ZN(new_n585_));
  OAI221_X1 g384(.A(new_n572_), .B1(new_n585_), .B2(new_n411_), .C1(new_n204_), .C2(new_n570_), .ZN(G1324gat));
  NOR2_X1   g385(.A1(new_n522_), .A2(new_n569_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(new_n412_), .A3(new_n396_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n396_), .B(new_n584_), .C1(new_n579_), .C2(new_n581_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(G8gat), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n589_), .B2(G8gat), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n588_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT40), .B(new_n588_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1325gat));
  NAND3_X1  g396(.A1(new_n587_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n582_), .A2(new_n244_), .A3(new_n584_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n599_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT41), .B1(new_n599_), .B2(G15gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(G1326gat));
  INV_X1    g401(.A(G22gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n587_), .A2(new_n603_), .A3(new_n397_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n582_), .A2(new_n397_), .A3(new_n584_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT42), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n605_), .A2(new_n606_), .A3(G22gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n605_), .B2(G22gat), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(G1327gat));
  NAND2_X1  g408(.A1(new_n552_), .A2(new_n567_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n520_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n436_), .A2(new_n611_), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n612_), .A2(G29gat), .A3(new_n372_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n521_), .A2(new_n567_), .A3(new_n434_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT103), .ZN(new_n615_));
  INV_X1    g414(.A(new_n553_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT43), .B1(new_n400_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n618_), .B(new_n553_), .C1(new_n395_), .C2(new_n399_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n615_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n373_), .B1(new_n620_), .B2(KEYINPUT44), .ZN(new_n621_));
  INV_X1    g420(.A(new_n615_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n618_), .B1(new_n577_), .B2(new_n553_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n619_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n622_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT104), .B(G29gat), .C1(new_n621_), .C2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n620_), .A2(KEYINPUT44), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n373_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT104), .B1(new_n632_), .B2(G29gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n613_), .B1(new_n629_), .B2(new_n633_), .ZN(G1328gat));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(KEYINPUT46), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n574_), .A2(G36gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n612_), .A2(KEYINPUT45), .A3(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT45), .B1(new_n612_), .B2(new_n638_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n574_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(new_n631_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n636_), .B1(new_n642_), .B2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n396_), .B1(new_n620_), .B2(KEYINPUT44), .ZN(new_n647_));
  OAI21_X1  g446(.A(G36gat), .B1(new_n647_), .B2(new_n627_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n641_), .C1(new_n635_), .C2(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1329gat));
  INV_X1    g449(.A(new_n244_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n232_), .B1(new_n612_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n630_), .A2(G43gat), .A3(new_n244_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n627_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT47), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT47), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n652_), .C1(new_n653_), .C2(new_n627_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1330gat));
  NAND3_X1  g457(.A1(new_n630_), .A2(new_n631_), .A3(new_n397_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n630_), .A2(new_n631_), .A3(KEYINPUT106), .A4(new_n397_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(G50gat), .A3(new_n662_), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n612_), .A2(G50gat), .A3(new_n355_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1331gat));
  NOR4_X1   g464(.A1(new_n569_), .A2(new_n400_), .A3(new_n521_), .A4(new_n434_), .ZN(new_n666_));
  INV_X1    g465(.A(G57gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n373_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n520_), .A2(new_n566_), .A3(new_n435_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n582_), .A2(new_n373_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n670_), .B2(new_n667_), .ZN(G1332gat));
  INV_X1    g470(.A(G64gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n672_), .A3(new_n396_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n582_), .A2(new_n396_), .A3(new_n669_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(G64gat), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G64gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1333gat));
  INV_X1    g477(.A(G71gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n666_), .A2(new_n679_), .A3(new_n244_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n582_), .A2(new_n244_), .A3(new_n669_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT49), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G71gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G71gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1334gat));
  NAND3_X1  g484(.A1(new_n666_), .A2(new_n349_), .A3(new_n397_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n582_), .A2(new_n397_), .A3(new_n669_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT50), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n687_), .A2(new_n688_), .A3(G78gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n687_), .B2(G78gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(G1335gat));
  NOR2_X1   g490(.A1(new_n400_), .A2(new_n434_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n610_), .A2(new_n521_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n455_), .A3(new_n373_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n567_), .A2(new_n520_), .A3(new_n583_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n373_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(new_n455_), .ZN(G1336gat));
  AOI21_X1  g499(.A(G92gat), .B1(new_n695_), .B2(new_n396_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n396_), .A2(G92gat), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT108), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n698_), .B2(new_n703_), .ZN(G1337gat));
  NAND3_X1  g503(.A1(new_n244_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n694_), .A2(new_n705_), .B1(KEYINPUT109), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n698_), .A2(new_n244_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G99gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(KEYINPUT109), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n709_), .B(new_n710_), .Z(G1338gat));
  AOI21_X1  g510(.A(new_n351_), .B1(KEYINPUT110), .B2(KEYINPUT52), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n698_), .B2(new_n397_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT53), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n716_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n695_), .A2(new_n351_), .A3(new_n397_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .A4(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n713_), .B(new_n715_), .C1(new_n698_), .C2(new_n397_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT53), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1339gat));
  AND4_X1   g524(.A1(new_n566_), .A2(new_n518_), .A3(new_n519_), .A4(new_n435_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n548_), .B(new_n726_), .C1(new_n552_), .C2(KEYINPUT37), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT54), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n432_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n424_), .A2(new_n419_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n423_), .B2(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n433_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n515_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT113), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n503_), .A2(new_n505_), .A3(new_n485_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n507_), .A2(KEYINPUT55), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n503_), .A2(new_n740_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n741_));
  AOI221_X4 g540(.A(new_n737_), .B1(new_n738_), .B2(new_n490_), .C1(new_n739_), .C2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n741_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n738_), .A2(new_n490_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT111), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n512_), .B1(new_n742_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n736_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT56), .B(new_n512_), .C1(new_n742_), .C2(new_n745_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n746_), .A2(new_n736_), .A3(new_n747_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n735_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT58), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT58), .B(new_n735_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n553_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n516_), .A2(new_n733_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n746_), .A2(new_n760_), .A3(new_n747_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n749_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n515_), .A2(new_n434_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n758_), .B1(new_n766_), .B2(new_n552_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n757_), .A2(new_n767_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n746_), .A2(new_n747_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT112), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n746_), .A2(new_n760_), .A3(new_n747_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n764_), .B1(new_n773_), .B2(new_n749_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT57), .B(new_n578_), .C1(new_n774_), .C2(new_n759_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n729_), .B1(new_n777_), .B2(new_n567_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n576_), .A2(new_n372_), .A3(new_n651_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n757_), .A2(new_n767_), .A3(new_n775_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n567_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n729_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n779_), .ZN(new_n786_));
  OAI22_X1  g585(.A1(new_n778_), .A2(new_n781_), .B1(new_n780_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G113gat), .B1(new_n787_), .B2(new_n435_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n434_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1340gat));
  OAI21_X1  g590(.A(G120gat), .B1(new_n787_), .B2(new_n521_), .ZN(new_n792_));
  INV_X1    g591(.A(G120gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n521_), .B2(KEYINPUT60), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n786_), .B(new_n794_), .C1(KEYINPUT60), .C2(new_n793_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n795_), .ZN(G1341gat));
  OAI21_X1  g595(.A(G127gat), .B1(new_n787_), .B2(new_n567_), .ZN(new_n797_));
  INV_X1    g596(.A(G127gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n786_), .A2(new_n798_), .A3(new_n566_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1342gat));
  AOI21_X1  g599(.A(G134gat), .B1(new_n786_), .B2(new_n552_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n787_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n553_), .A2(G134gat), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT116), .Z(new_n804_));
  AOI21_X1  g603(.A(new_n801_), .B1(new_n802_), .B2(new_n804_), .ZN(G1343gat));
  NAND4_X1  g604(.A1(new_n574_), .A2(new_n373_), .A3(new_n397_), .A4(new_n651_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT117), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n785_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n434_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n808_), .B2(new_n520_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n785_), .A2(new_n807_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n813_), .A2(KEYINPUT119), .A3(new_n521_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT118), .B(G148gat), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OR3_X1    g615(.A1(new_n812_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1345gat));
  NOR2_X1   g618(.A1(new_n813_), .A2(new_n567_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT61), .B(G155gat), .Z(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1346gat));
  AOI21_X1  g621(.A(G162gat), .B1(new_n808_), .B2(new_n552_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n553_), .A2(G162gat), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT120), .Z(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n808_), .B2(new_n825_), .ZN(G1347gat));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n212_), .B1(new_n827_), .B2(KEYINPUT62), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n574_), .A2(new_n398_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n397_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n434_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n778_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(KEYINPUT121), .A3(new_n834_), .ZN(new_n835_));
  OAI221_X1 g634(.A(new_n828_), .B1(new_n827_), .B2(KEYINPUT62), .C1(new_n778_), .C2(new_n832_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n778_), .A2(new_n832_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n227_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n836_), .A3(new_n838_), .ZN(G1348gat));
  INV_X1    g638(.A(new_n831_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n778_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n520_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n729_), .B1(new_n782_), .B2(new_n567_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n397_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n830_), .A2(new_n213_), .A3(new_n521_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n842_), .A2(new_n226_), .B1(new_n844_), .B2(new_n845_), .ZN(G1349gat));
  NOR2_X1   g645(.A1(new_n830_), .A2(new_n567_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G183gat), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n567_), .A2(new_n205_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n841_), .B2(new_n849_), .ZN(G1350gat));
  NAND3_X1  g649(.A1(new_n841_), .A2(new_n206_), .A3(new_n552_), .ZN(new_n851_));
  INV_X1    g650(.A(G190gat), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n778_), .A2(new_n616_), .A3(new_n840_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1351gat));
  NAND3_X1  g653(.A1(new_n396_), .A2(new_n374_), .A3(new_n651_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT122), .B1(new_n785_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n843_), .A2(new_n858_), .A3(new_n855_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT123), .B(new_n261_), .C1(new_n860_), .C2(new_n583_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n785_), .A2(KEYINPUT122), .A3(new_n856_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n858_), .B1(new_n843_), .B2(new_n855_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n583_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G197gat), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n864_), .B2(G197gat), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n861_), .A2(new_n865_), .A3(new_n867_), .ZN(G1352gat));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n863_), .ZN(new_n869_));
  INV_X1    g668(.A(G204gat), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n869_), .B(new_n520_), .C1(KEYINPUT124), .C2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n860_), .A2(new_n521_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT124), .B(G204gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1353gat));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  NAND2_X1  g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n566_), .A2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT125), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n869_), .B2(new_n881_), .ZN(new_n882_));
  AOI211_X1 g681(.A(KEYINPUT126), .B(new_n880_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n876_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n881_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT126), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n869_), .A2(new_n877_), .A3(new_n881_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n875_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n888_), .ZN(G1354gat));
  AOI21_X1  g688(.A(G218gat), .B1(new_n869_), .B2(new_n552_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n553_), .A2(G218gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT127), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n869_), .B2(new_n892_), .ZN(G1355gat));
endmodule


