//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT11), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n206_));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n202_), .A3(KEYINPUT11), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .A4(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(KEYINPUT11), .B2(new_n203_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(new_n204_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  OAI22_X1  g012(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n214_), .B(new_n217_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n220_), .B(KEYINPUT6), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n225_), .A2(KEYINPUT67), .A3(new_n214_), .A4(new_n217_), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  INV_X1    g026(.A(G92gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n229_), .A2(KEYINPUT8), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n224_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n219_), .A2(new_n221_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n217_), .A2(new_n214_), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT68), .B(new_n233_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT8), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT68), .B1(new_n222_), .B2(new_n233_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n232_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(G85gat), .B2(G92gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n227_), .A2(KEYINPUT64), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G85gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT9), .B1(new_n245_), .B2(G92gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n241_), .B1(new_n246_), .B2(KEYINPUT65), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT64), .B(G85gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(new_n228_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n250_), .B2(KEYINPUT9), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT10), .B(G99gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n225_), .B1(G106gat), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n213_), .B1(new_n239_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT12), .B1(new_n257_), .B2(KEYINPUT71), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n254_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n222_), .A2(new_n233_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(KEYINPUT8), .A3(new_n236_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n265_), .B2(new_n232_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n259_), .B(new_n260_), .C1(new_n266_), .C2(new_n213_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n213_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n258_), .A2(new_n267_), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n257_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n239_), .A2(new_n256_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n213_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT70), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n272_), .B1(new_n257_), .B2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G176gat), .B(G204gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT73), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G120gat), .B(G148gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n270_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT74), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n270_), .A2(new_n276_), .A3(new_n285_), .A4(new_n282_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n270_), .A2(new_n276_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n282_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n287_), .A2(KEYINPUT13), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT13), .B1(new_n287_), .B2(new_n290_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G15gat), .B(G22gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT81), .B(G1gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT82), .B(G8gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n294_), .B1(new_n297_), .B2(KEYINPUT14), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G29gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G43gat), .B(G50gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT15), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n300_), .A2(new_n304_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G229gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT87), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT86), .B1(new_n300_), .B2(new_n304_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n304_), .B2(new_n300_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n304_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n301_), .A2(KEYINPUT86), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n306_), .A2(new_n317_), .A3(new_n309_), .A4(new_n307_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G113gat), .B(G141gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G169gat), .B(G197gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n311_), .A2(new_n316_), .A3(new_n318_), .A4(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n293_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT90), .B1(G169gat), .B2(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT24), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G183gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT25), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(KEYINPUT25), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G190gat), .ZN(new_n340_));
  OR3_X1    g139(.A1(new_n340_), .A2(KEYINPUT89), .A3(KEYINPUT26), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(new_n342_), .A3(G183gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT26), .B1(new_n340_), .B2(KEYINPUT89), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n334_), .B1(new_n339_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT91), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT23), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n330_), .A2(new_n350_), .A3(new_n331_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n346_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n347_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n349_), .B1(G183gat), .B2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(G176gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(KEYINPUT92), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G169gat), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(G169gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n355_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT93), .B(G43gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n363_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(G15gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT30), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(KEYINPUT94), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT94), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT101), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G22gat), .B(G50gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G141gat), .A2(G148gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT95), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G141gat), .A2(G148gat), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT1), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(G155gat), .A3(G162gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT97), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(G155gat), .B2(G162gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT96), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(KEYINPUT96), .A3(new_n400_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n394_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT98), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n393_), .B(KEYINPUT3), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n407_), .B(new_n408_), .C1(KEYINPUT2), .C2(new_n392_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G155gat), .B(G162gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT99), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n404_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n416_), .A2(KEYINPUT28), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(KEYINPUT28), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n390_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n416_), .A2(KEYINPUT28), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(KEYINPUT28), .ZN(new_n421_));
  INV_X1    g220(.A(new_n390_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n389_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G197gat), .B(G204gat), .Z(new_n426_));
  OR2_X1    g225(.A1(new_n426_), .A2(KEYINPUT21), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(KEYINPUT21), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G211gat), .B(G218gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n428_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT100), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT29), .B1(new_n404_), .B2(new_n413_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n432_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n435_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n388_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n419_), .A2(new_n423_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n425_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n441_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n419_), .A2(new_n423_), .A3(new_n442_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n424_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT104), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT103), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n414_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n371_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n414_), .A2(new_n453_), .A3(new_n370_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n414_), .A2(KEYINPUT4), .A3(new_n371_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(new_n450_), .A3(new_n456_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G85gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT0), .B(G57gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n449_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n459_), .A2(new_n460_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n464_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT104), .A3(new_n466_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n448_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT102), .ZN(new_n476_));
  INV_X1    g275(.A(new_n337_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n477_), .A2(new_n336_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT26), .B(G190gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n480_), .A2(new_n334_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n481_), .A2(new_n352_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n333_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT22), .B(G169gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n357_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n356_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n476_), .B(new_n432_), .C1(new_n482_), .C2(new_n486_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n481_), .A2(new_n352_), .B1(new_n356_), .B2(new_n485_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n432_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT102), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n432_), .B(KEYINPUT100), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT20), .B1(new_n493_), .B2(new_n363_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n475_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G8gat), .B(G36gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT18), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G64gat), .B(G92gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n363_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n434_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n495_), .B(new_n499_), .C1(new_n475_), .C2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n499_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n475_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n500_), .B1(new_n502_), .B2(new_n434_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(new_n491_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n503_), .A2(new_n475_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT27), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n507_), .A2(new_n506_), .A3(new_n491_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n503_), .A2(new_n475_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n505_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n504_), .A3(KEYINPUT27), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n473_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n455_), .A2(new_n456_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT4), .ZN(new_n522_));
  INV_X1    g321(.A(new_n458_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n450_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n464_), .B1(new_n521_), .B2(new_n451_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n504_), .A2(new_n510_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT33), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n471_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n468_), .A2(KEYINPUT33), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n516_), .A2(KEYINPUT32), .A3(new_n499_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n499_), .A2(KEYINPUT32), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n495_), .B(new_n533_), .C1(new_n475_), .C2(new_n503_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(new_n534_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n448_), .B1(new_n531_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n387_), .B1(new_n520_), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n519_), .A2(new_n448_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n469_), .A2(new_n472_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n540_), .A3(new_n383_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n327_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n239_), .A2(new_n256_), .A3(new_n304_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(KEYINPUT34), .Z(new_n545_));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT75), .Z(new_n548_));
  INV_X1    g347(.A(new_n305_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n543_), .B(new_n548_), .C1(new_n266_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT77), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT76), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n273_), .A2(new_n305_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT76), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n543_), .A4(new_n548_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n545_), .A2(new_n546_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  OAI221_X1 g356(.A(KEYINPUT76), .B1(new_n546_), .B2(new_n545_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT78), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(KEYINPUT78), .A3(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n562_), .B(KEYINPUT36), .Z(new_n569_));
  NAND3_X1  g368(.A1(new_n557_), .A2(new_n569_), .A3(new_n558_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(KEYINPUT37), .A3(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n557_), .A2(KEYINPUT79), .A3(new_n558_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT79), .B1(new_n557_), .B2(new_n558_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n569_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT80), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(KEYINPUT80), .B(new_n569_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(new_n568_), .A3(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n571_), .B1(new_n578_), .B2(KEYINPUT37), .ZN(new_n579_));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT17), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT85), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(new_n213_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n301_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT83), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n584_), .A2(KEYINPUT17), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n579_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n542_), .A2(new_n596_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n597_), .A2(new_n295_), .A3(new_n540_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT38), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT106), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n578_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n594_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT105), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n327_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT105), .B1(new_n293_), .B2(new_n326_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n539_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n599_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n601_), .A2(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n519_), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n597_), .A2(new_n296_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n519_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(KEYINPUT107), .A2(KEYINPUT39), .ZN(new_n615_));
  INV_X1    g414(.A(G8gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(KEYINPUT107), .B2(KEYINPUT39), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n614_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n615_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(G1325gat));
  INV_X1    g421(.A(new_n387_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n376_), .B1(new_n608_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT41), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n376_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n597_), .B2(new_n626_), .ZN(G1326gat));
  INV_X1    g426(.A(G22gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n608_), .B2(new_n448_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT42), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n448_), .A2(new_n628_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT108), .Z(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n597_), .B2(new_n632_), .ZN(G1327gat));
  NAND3_X1  g432(.A1(new_n576_), .A2(new_n568_), .A3(new_n577_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n594_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n542_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n539_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n537_), .A2(new_n541_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n579_), .ZN(new_n640_));
  XOR2_X1   g439(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n639_), .B(new_n579_), .C1(KEYINPUT109), .C2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n595_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT44), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n649_), .B(new_n646_), .C1(new_n642_), .C2(new_n644_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(KEYINPUT110), .A3(new_n539_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT110), .B1(new_n651_), .B2(new_n539_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n638_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(G36gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n636_), .A2(new_n656_), .A3(new_n519_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n648_), .A2(new_n650_), .A3(new_n612_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n656_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n658_), .B(KEYINPUT46), .C1(new_n659_), .C2(new_n656_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  INV_X1    g463(.A(KEYINPUT47), .ZN(new_n665_));
  INV_X1    g464(.A(G43gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n651_), .B2(new_n383_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n636_), .A2(new_n666_), .A3(new_n623_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n645_), .A2(new_n647_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n649_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n645_), .A2(KEYINPUT44), .A3(new_n647_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n383_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G43gat), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(KEYINPUT47), .A3(new_n668_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n670_), .A2(new_n677_), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n636_), .B2(new_n448_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n448_), .A2(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n651_), .B2(new_n680_), .ZN(G1331gat));
  NOR2_X1   g480(.A1(new_n293_), .A2(new_n326_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n639_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n596_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n539_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT111), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n602_), .A2(new_n594_), .A3(new_n682_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(G57gat), .A3(new_n539_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1332gat));
  INV_X1    g488(.A(G64gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n687_), .B2(new_n519_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n690_), .A3(new_n519_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1333gat));
  INV_X1    g494(.A(G71gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n687_), .B2(new_n623_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT49), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n684_), .A2(new_n696_), .A3(new_n623_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1334gat));
  INV_X1    g499(.A(G78gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n687_), .B2(new_n448_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT50), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n684_), .A2(new_n701_), .A3(new_n448_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1335gat));
  NAND2_X1  g504(.A1(new_n683_), .A2(new_n635_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n227_), .B1(new_n706_), .B2(new_n540_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT113), .Z(new_n708_));
  NAND2_X1  g507(.A1(new_n682_), .A2(new_n595_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT114), .Z(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n712_), .A2(new_n249_), .A3(new_n540_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n708_), .A2(new_n713_), .ZN(G1336gat));
  OAI21_X1  g513(.A(new_n228_), .B1(new_n706_), .B2(new_n612_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT115), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n712_), .A2(new_n228_), .A3(new_n612_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1337gat));
  NOR3_X1   g517(.A1(new_n706_), .A2(new_n253_), .A3(new_n675_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n711_), .A2(new_n623_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G99gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(G1338gat));
  INV_X1    g522(.A(G106gat), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n683_), .A2(new_n724_), .A3(new_n448_), .A4(new_n635_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n711_), .A2(new_n448_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G106gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT52), .B(new_n724_), .C1(new_n711_), .C2(new_n448_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT53), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT53), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(new_n725_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1339gat));
  NAND3_X1  g533(.A1(new_n538_), .A2(new_n539_), .A3(new_n383_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(KEYINPUT59), .ZN(new_n736_));
  INV_X1    g535(.A(new_n569_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT79), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n559_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n557_), .A2(KEYINPUT79), .A3(new_n558_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n741_), .A2(KEYINPUT80), .B1(new_n566_), .B2(new_n567_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT37), .B1(new_n742_), .B2(new_n576_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n571_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n326_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n745_), .A2(new_n594_), .A3(new_n746_), .A4(new_n293_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n747_), .B(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n287_), .A2(new_n326_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n258_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n268_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n270_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n753_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n289_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n273_), .A2(new_n274_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n259_), .B1(new_n266_), .B2(new_n213_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(KEYINPUT12), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n268_), .B1(new_n764_), .B2(new_n267_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n270_), .B1(new_n765_), .B2(new_n752_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n758_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n289_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n751_), .B1(new_n761_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n313_), .A2(new_n309_), .A3(new_n315_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n323_), .C1(new_n309_), .C2(new_n308_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n325_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n567_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT78), .B1(new_n559_), .B2(new_n563_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n577_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n741_), .A2(KEYINPUT80), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n770_), .A2(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n773_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n287_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n287_), .A2(new_n782_), .A3(KEYINPUT120), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n768_), .B2(new_n289_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n760_), .B(new_n282_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n785_), .B(new_n786_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n761_), .A2(new_n769_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n791_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n792_), .B(new_n795_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n781_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n751_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n774_), .B1(new_n793_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT118), .B1(new_n799_), .B2(new_n578_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n634_), .B(new_n801_), .C1(new_n770_), .C2(new_n774_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n780_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n594_), .B1(new_n797_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n736_), .B1(new_n750_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n796_), .A2(KEYINPUT122), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT122), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n579_), .A2(new_n807_), .A3(new_n795_), .A4(new_n792_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n803_), .A2(KEYINPUT119), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT57), .B1(new_n779_), .B2(KEYINPUT118), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n802_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n809_), .A2(new_n810_), .A3(new_n781_), .A4(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n595_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n750_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n735_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n805_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n746_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n816_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n735_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OR3_X1    g622(.A1(new_n823_), .A2(G113gat), .A3(new_n746_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n820_), .A2(new_n824_), .ZN(G1340gat));
  XOR2_X1   g624(.A(KEYINPUT123), .B(G120gat), .Z(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n293_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n817_), .B(new_n827_), .C1(KEYINPUT60), .C2(new_n826_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n819_), .A2(new_n293_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n826_), .ZN(G1341gat));
  OAI21_X1  g629(.A(G127gat), .B1(new_n819_), .B2(new_n595_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n823_), .A2(G127gat), .A3(new_n595_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1342gat));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n634_), .B(new_n735_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G134gat), .ZN(new_n836_));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT124), .B(new_n837_), .C1(new_n823_), .C2(new_n634_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n750_), .A2(new_n804_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n823_), .A2(KEYINPUT59), .B1(new_n839_), .B2(new_n736_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n745_), .A2(new_n837_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n836_), .A2(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(G1343gat));
  AND4_X1   g641(.A1(new_n448_), .A2(new_n387_), .A3(new_n539_), .A4(new_n612_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n821_), .A2(new_n326_), .A3(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g644(.A(new_n293_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n821_), .A2(new_n846_), .A3(new_n843_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT125), .B(G148gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n847_), .B(new_n848_), .Z(G1345gat));
  AND4_X1   g648(.A1(new_n812_), .A2(new_n800_), .A3(new_n780_), .A4(new_n802_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n812_), .B1(new_n811_), .B2(new_n802_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n781_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n594_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n594_), .B(new_n843_), .C1(new_n855_), .C2(new_n750_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT126), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT126), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n821_), .A2(new_n858_), .A3(new_n594_), .A4(new_n843_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n857_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1346gat));
  NAND2_X1  g662(.A1(new_n821_), .A2(new_n843_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G162gat), .B1(new_n864_), .B2(new_n745_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n634_), .A2(G162gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n864_), .B2(new_n866_), .ZN(G1347gat));
  NAND3_X1  g666(.A1(new_n623_), .A2(new_n540_), .A3(new_n519_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT127), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n448_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n839_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G169gat), .B1(new_n871_), .B2(new_n746_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n839_), .A2(new_n870_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n326_), .A3(new_n484_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT62), .B(G169gat), .C1(new_n871_), .C2(new_n746_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n875_), .B2(new_n846_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n448_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n869_), .A2(new_n357_), .A3(new_n293_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(G1349gat));
  NOR3_X1   g681(.A1(new_n871_), .A2(new_n595_), .A3(new_n478_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n869_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n594_), .A3(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n335_), .B2(new_n885_), .ZN(G1350gat));
  NAND3_X1  g685(.A1(new_n875_), .A2(new_n578_), .A3(new_n479_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G190gat), .B1(new_n871_), .B2(new_n745_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n623_), .A2(new_n473_), .A3(new_n612_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n821_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G197gat), .B1(new_n892_), .B2(new_n326_), .ZN(new_n893_));
  INV_X1    g692(.A(G197gat), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n891_), .A2(new_n894_), .A3(new_n746_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1352gat));
  OR3_X1    g695(.A1(new_n891_), .A2(G204gat), .A3(new_n293_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G204gat), .B1(new_n891_), .B2(new_n293_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1353gat));
  XNOR2_X1  g698(.A(KEYINPUT63), .B(G211gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n891_), .A2(new_n595_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n892_), .A2(new_n594_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1354gat));
  OR3_X1    g703(.A1(new_n891_), .A2(G218gat), .A3(new_n634_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G218gat), .B1(new_n891_), .B2(new_n745_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1355gat));
endmodule


