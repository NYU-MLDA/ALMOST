//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G85gat), .Z(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n212_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT10), .B(G99gat), .Z(new_n220_));
  AOI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT66), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT7), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n212_), .A2(new_n214_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(KEYINPUT8), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n223_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n230_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n222_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n207_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n206_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT34), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT68), .B(KEYINPUT35), .Z(new_n242_));
  OAI211_X1 g041(.A(new_n237_), .B(new_n239_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(KEYINPUT69), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(new_n245_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G190gat), .B(G218gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G134gat), .ZN(new_n250_));
  INV_X1    g049(.A(G162gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI22_X1  g052(.A1(new_n247_), .A2(new_n248_), .B1(KEYINPUT36), .B2(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n243_), .A2(new_n245_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n252_), .B(KEYINPUT36), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n257_), .A3(new_n246_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT37), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT37), .ZN(new_n262_));
  AOI211_X1 g061(.A(KEYINPUT70), .B(new_n262_), .C1(new_n254_), .C2(new_n258_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT11), .ZN(new_n266_));
  XOR2_X1   g065(.A(G71gat), .B(G78gat), .Z(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n265_), .A2(KEYINPUT11), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n269_), .A2(new_n266_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n270_), .B2(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G231gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G1gat), .B(G8gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT71), .ZN(new_n275_));
  INV_X1    g074(.A(G15gat), .ZN(new_n276_));
  INV_X1    g075(.A(G22gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G15gat), .A2(G22gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G1gat), .A2(G8gat), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n278_), .A2(new_n279_), .B1(KEYINPUT14), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n275_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n273_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G127gat), .B(G155gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G183gat), .B(G211gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT17), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n283_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n288_), .B(new_n289_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n283_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT73), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n264_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT74), .Z(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(G113gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(G113gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n299_), .A2(G120gat), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(G120gat), .B1(new_n299_), .B2(new_n300_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT31), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT79), .B(G176gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT22), .B(G169gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(KEYINPUT23), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(KEYINPUT23), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n312_), .B1(new_n316_), .B2(new_n310_), .ZN(new_n317_));
  AND2_X1   g116(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n318_), .A2(new_n319_), .A3(G190gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n309_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT76), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n323_), .B(KEYINPUT25), .C1(KEYINPUT76), .C2(G183gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(KEYINPUT24), .A3(new_n305_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n313_), .A2(new_n315_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n329_), .A2(KEYINPUT78), .A3(KEYINPUT24), .A4(new_n305_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n328_), .A2(new_n332_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n321_), .A2(new_n322_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n322_), .B1(new_n321_), .B2(new_n337_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G15gat), .B(G43gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G99gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G71gat), .ZN(new_n344_));
  INV_X1    g143(.A(G71gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G99gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n344_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n342_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n346_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n347_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n344_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n341_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n340_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n350_), .A2(new_n355_), .A3(new_n340_), .ZN(new_n357_));
  OAI22_X1  g156(.A1(new_n338_), .A2(new_n339_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n321_), .A2(new_n337_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT30), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n321_), .A2(new_n322_), .A3(new_n337_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n358_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n304_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT84), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(new_n363_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n369_), .A2(new_n304_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n371_), .B(new_n304_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT85), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n368_), .A2(new_n375_), .A3(new_n370_), .A4(new_n372_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT95), .ZN(new_n378_));
  OR2_X1    g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT86), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G141gat), .A3(G148gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G141gat), .ZN(new_n388_));
  INV_X1    g187(.A(G148gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n387_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT2), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT89), .B1(new_n383_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT89), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n395_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398_));
  OAI22_X1  g197(.A1(new_n398_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(KEYINPUT87), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n398_), .A2(new_n388_), .A3(new_n389_), .A4(KEYINPUT3), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n397_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT88), .B1(new_n387_), .B2(new_n393_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407_));
  AOI211_X1 g206(.A(new_n407_), .B(KEYINPUT2), .C1(new_n384_), .C2(new_n386_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n405_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n379_), .A2(new_n381_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n378_), .B(new_n392_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n303_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n392_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n387_), .A2(new_n393_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n407_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n387_), .A2(KEYINPUT88), .A3(new_n393_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n398_), .A2(KEYINPUT3), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n400_), .A2(KEYINPUT87), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n390_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n420_), .A2(new_n403_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n416_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n410_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n414_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n378_), .A3(new_n303_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n413_), .A2(KEYINPUT4), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT96), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n424_), .A2(KEYINPUT4), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(new_n412_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n413_), .A2(new_n427_), .A3(new_n425_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT0), .B(G57gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G85gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(G1gat), .B(G29gat), .Z(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n377_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT29), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n424_), .B2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n406_), .A2(new_n408_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n410_), .B1(new_n445_), .B2(new_n421_), .ZN(new_n446_));
  OAI211_X1 g245(.A(KEYINPUT91), .B(KEYINPUT29), .C1(new_n446_), .C2(new_n414_), .ZN(new_n447_));
  INV_X1    g246(.A(G204gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G197gat), .ZN(new_n449_));
  INV_X1    g248(.A(G197gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G204gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT21), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT21), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n449_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G211gat), .B(G218gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G211gat), .B(G218gat), .Z(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT21), .A3(new_n452_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n444_), .A2(new_n447_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G228gat), .ZN(new_n462_));
  INV_X1    g261(.A(G233gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n424_), .A2(new_n443_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n457_), .A2(KEYINPUT90), .A3(new_n459_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT90), .B1(new_n457_), .B2(new_n459_), .ZN(new_n469_));
  OAI22_X1  g268(.A1(new_n468_), .A2(new_n469_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n465_), .A2(KEYINPUT92), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G78gat), .B(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n465_), .A2(new_n472_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT92), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n443_), .B(new_n392_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT28), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT28), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n424_), .A2(new_n481_), .A3(new_n443_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G22gat), .B(G50gat), .Z(new_n483_));
  AND3_X1   g282(.A1(new_n480_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n471_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n474_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT92), .A3(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n475_), .A2(new_n478_), .A3(new_n486_), .A4(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n486_), .B1(KEYINPUT92), .B2(new_n487_), .ZN(new_n491_));
  AND4_X1   g290(.A1(KEYINPUT92), .A2(new_n465_), .A3(new_n472_), .A4(new_n488_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n488_), .B1(new_n487_), .B2(KEYINPUT92), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n455_), .A2(new_n456_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n454_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n458_), .A2(KEYINPUT21), .A3(new_n452_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n496_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n501_), .A2(new_n321_), .A3(new_n337_), .A4(new_n467_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT19), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(KEYINPUT24), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n334_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(KEYINPUT24), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n329_), .A2(new_n510_), .A3(new_n511_), .A4(new_n305_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n325_), .A2(G183gat), .ZN(new_n513_));
  INV_X1    g312(.A(G183gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT25), .ZN(new_n515_));
  AND2_X1   g314(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n513_), .B(new_n515_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n509_), .A2(new_n512_), .A3(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT79), .B(G176gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n305_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G183gat), .A2(G190gat), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n526_));
  OAI22_X1  g325(.A1(new_n519_), .A2(new_n317_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n460_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n502_), .A2(KEYINPUT20), .A3(new_n505_), .A4(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT20), .B1(new_n527_), .B2(new_n460_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n360_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n534_));
  OAI211_X1 g333(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n527_), .C2(new_n460_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n530_), .B1(new_n504_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT18), .B(G64gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G92gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G8gat), .B(G36gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT27), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n502_), .A2(KEYINPUT20), .A3(new_n528_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n504_), .ZN(new_n544_));
  OAI211_X1 g343(.A(KEYINPUT20), .B(new_n505_), .C1(new_n527_), .C2(new_n460_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n534_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n544_), .A2(new_n541_), .A3(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT99), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT27), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n536_), .A2(new_n504_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n529_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n541_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT99), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n543_), .A2(new_n504_), .B1(new_n546_), .B2(new_n534_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n541_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n549_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n556_), .B2(new_n541_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n544_), .A2(new_n547_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n553_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n560_), .A3(new_n553_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n495_), .A2(new_n559_), .A3(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n441_), .A2(new_n568_), .A3(KEYINPUT101), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT101), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n490_), .A2(new_n494_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n555_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n541_), .B1(new_n551_), .B2(new_n529_), .ZN(new_n573_));
  NOR4_X1   g372(.A1(new_n573_), .A2(new_n548_), .A3(KEYINPUT99), .A4(new_n550_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n567_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n440_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n570_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n575_), .A2(new_n495_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n541_), .A2(KEYINPUT32), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n556_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n537_), .B2(new_n582_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n440_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n564_), .A2(new_n565_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n429_), .A2(new_n412_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n426_), .A2(new_n427_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n413_), .A2(new_n425_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n588_), .B(new_n436_), .C1(new_n589_), .C2(new_n428_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n431_), .A2(KEYINPUT33), .A3(new_n432_), .A4(new_n437_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n586_), .A2(new_n590_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n583_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n582_), .B1(new_n551_), .B2(new_n529_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n598_), .B(KEYINPUT98), .C1(new_n439_), .C2(new_n438_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n585_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n580_), .A2(new_n440_), .B1(new_n600_), .B2(new_n495_), .ZN(new_n601_));
  OAI22_X1  g400(.A1(new_n569_), .A2(new_n579_), .B1(new_n601_), .B2(new_n377_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n236_), .A2(KEYINPUT12), .A3(new_n271_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(G230gat), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n236_), .A2(new_n271_), .B1(new_n605_), .B2(new_n463_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT12), .B1(new_n236_), .B2(new_n271_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n604_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n605_), .A2(new_n463_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n236_), .A2(new_n271_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n236_), .A2(new_n271_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n448_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(G176gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT67), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n615_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT13), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n207_), .A2(new_n282_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n238_), .A2(new_n282_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n238_), .B(new_n282_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(G229gat), .A3(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G113gat), .B(G141gat), .ZN(new_n629_));
  INV_X1    g428(.A(G169gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n450_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n626_), .A2(new_n628_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT75), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n626_), .A2(new_n628_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n632_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n635_), .B(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n622_), .A2(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n602_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n297_), .A2(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n642_), .A2(G1gat), .A3(new_n440_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n643_), .A2(KEYINPUT38), .ZN(new_n644_));
  INV_X1    g443(.A(new_n259_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n602_), .A2(new_n645_), .A3(new_n640_), .A4(new_n294_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n440_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(KEYINPUT38), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT102), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n644_), .A2(new_n651_), .A3(new_n647_), .A4(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1324gat));
  AND2_X1   g452(.A1(new_n564_), .A2(new_n565_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n549_), .A2(new_n558_), .B1(new_n654_), .B2(new_n566_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n642_), .A2(G8gat), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G8gat), .B1(new_n646_), .B2(new_n655_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g460(.A(new_n377_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G15gat), .B1(new_n646_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  INV_X1    g463(.A(new_n642_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n276_), .A3(new_n377_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1326gat));
  XNOR2_X1  g466(.A(new_n495_), .B(KEYINPUT103), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n277_), .A3(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n646_), .A2(new_n668_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G22gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT104), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n674_), .A3(G22gat), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n673_), .A2(KEYINPUT42), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT42), .B1(new_n673_), .B2(new_n675_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n670_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT105), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n670_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1327gat));
  NOR3_X1   g481(.A1(new_n622_), .A2(new_n639_), .A3(new_n295_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT106), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT106), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n600_), .A2(new_n495_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n655_), .A2(new_n571_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n577_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n662_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT101), .B1(new_n441_), .B2(new_n568_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n576_), .A2(new_n570_), .A3(new_n578_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT43), .B(new_n264_), .C1(new_n690_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n261_), .A2(new_n263_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n602_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n686_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n686_), .C1(new_n694_), .C2(new_n697_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n577_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n700_), .A2(KEYINPUT107), .A3(new_n577_), .A4(new_n701_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(G29gat), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(G29gat), .A4(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n295_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n259_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT109), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n641_), .A2(new_n713_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n714_), .A2(G29gat), .A3(new_n440_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n710_), .A2(new_n715_), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n714_), .A2(G36gat), .A3(new_n655_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n700_), .A2(new_n701_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n655_), .ZN(new_n721_));
  INV_X1    g520(.A(G36gat), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n719_), .B(KEYINPUT46), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n721_), .A2(new_n722_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n718_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1329gat));
  NOR3_X1   g526(.A1(new_n714_), .A2(G43gat), .A3(new_n662_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n700_), .A2(new_n377_), .A3(new_n701_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G43gat), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n720_), .B2(new_n495_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n669_), .A2(new_n205_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n714_), .B2(new_n733_), .ZN(G1331gat));
  NAND2_X1  g533(.A1(new_n297_), .A2(new_n622_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n735_), .A2(KEYINPUT110), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n638_), .B1(new_n735_), .B2(KEYINPUT110), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n602_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n577_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n622_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n638_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n602_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n645_), .A3(new_n295_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n440_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n739_), .B1(G57gat), .B2(new_n744_), .ZN(G1332gat));
  INV_X1    g544(.A(G64gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n738_), .A2(new_n746_), .A3(new_n575_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G64gat), .B1(new_n743_), .B2(new_n655_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT48), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1333gat));
  NAND3_X1  g549(.A1(new_n738_), .A2(new_n345_), .A3(new_n377_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G71gat), .B1(new_n743_), .B2(new_n662_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT49), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1334gat));
  INV_X1    g553(.A(G78gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n738_), .A2(new_n755_), .A3(new_n669_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G78gat), .B1(new_n743_), .B2(new_n668_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1335gat));
  AND2_X1   g558(.A1(new_n742_), .A2(new_n713_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n577_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n694_), .A2(new_n697_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n762_), .A2(new_n711_), .A3(new_n741_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n440_), .A2(new_n209_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  NAND3_X1  g564(.A1(new_n763_), .A2(G92gat), .A3(new_n575_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n760_), .A2(new_n575_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(KEYINPUT111), .A3(new_n210_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT111), .B1(new_n767_), .B2(new_n210_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT112), .ZN(G1337gat));
  NAND4_X1  g570(.A1(new_n762_), .A2(new_n377_), .A3(new_n711_), .A4(new_n741_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n772_), .A2(KEYINPUT113), .A3(G99gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT113), .B1(new_n772_), .B2(G99gat), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(KEYINPUT114), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n760_), .A2(new_n220_), .A3(new_n377_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n772_), .A2(G99gat), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n772_), .A2(KEYINPUT113), .A3(G99gat), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .A4(new_n777_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n778_), .A2(new_n785_), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n760_), .A2(new_n219_), .A3(new_n571_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n762_), .A2(new_n571_), .A3(new_n711_), .A4(new_n741_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(G106gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n788_), .B2(G106gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n787_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  NOR3_X1   g595(.A1(new_n662_), .A2(new_n568_), .A3(new_n440_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n294_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n603_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(KEYINPUT55), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n610_), .A2(KEYINPUT116), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n604_), .A2(new_n609_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n611_), .B1(new_n806_), .B2(new_n613_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n802_), .A2(KEYINPUT55), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n803_), .A2(new_n805_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n619_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n619_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n627_), .A2(new_n624_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n623_), .A2(new_n625_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n632_), .B(new_n816_), .C1(new_n817_), .C2(new_n624_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n634_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n615_), .A2(new_n619_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n800_), .B1(new_n815_), .B2(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n821_), .B(KEYINPUT119), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT58), .A3(new_n814_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n696_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n619_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n820_), .B1(new_n828_), .B2(KEYINPUT117), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n638_), .B(new_n829_), .C1(new_n814_), .C2(KEYINPUT117), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n621_), .A2(new_n819_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n259_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n827_), .B1(new_n834_), .B2(KEYINPUT57), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n836_), .B(new_n259_), .C1(new_n830_), .C2(new_n833_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n799_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n639_), .A2(new_n295_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT115), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n696_), .A2(new_n840_), .A3(new_n622_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(KEYINPUT115), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n264_), .B(new_n740_), .C1(KEYINPUT115), .C2(new_n839_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n843_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n798_), .B1(new_n838_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849_), .B2(new_n638_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n835_), .A2(KEYINPUT120), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n827_), .B(new_n852_), .C1(new_n834_), .C2(KEYINPUT57), .ZN(new_n853_));
  INV_X1    g652(.A(new_n837_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n711_), .B1(new_n851_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n848_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n838_), .A2(new_n848_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n797_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n857_), .A2(new_n858_), .B1(new_n860_), .B2(KEYINPUT59), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n861_), .A2(G113gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n850_), .B1(new_n862_), .B2(new_n638_), .ZN(G1340gat));
  NAND2_X1  g662(.A1(new_n835_), .A2(KEYINPUT120), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n854_), .A3(new_n853_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n865_), .A2(new_n711_), .B1(new_n847_), .B2(new_n844_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n858_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n868_), .B2(new_n849_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G120gat), .B1(new_n869_), .B2(new_n740_), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n849_), .B1(KEYINPUT60), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n740_), .B2(KEYINPUT60), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT121), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n870_), .B1(new_n872_), .B2(new_n874_), .ZN(G1341gat));
  AOI21_X1  g674(.A(G127gat), .B1(new_n849_), .B2(new_n295_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n294_), .A2(G127gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n861_), .B2(new_n877_), .ZN(G1342gat));
  AOI21_X1  g677(.A(new_n867_), .B1(new_n856_), .B2(new_n848_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n849_), .A2(new_n868_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n696_), .A2(G134gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G134gat), .B1(new_n849_), .B2(new_n259_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  INV_X1    g684(.A(new_n883_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n885_), .B(new_n886_), .C1(new_n869_), .C2(new_n881_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(G1343gat));
  AOI21_X1  g687(.A(new_n377_), .B1(new_n838_), .B2(new_n848_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n639_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n388_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n740_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n389_), .ZN(G1345gat));
  NOR2_X1   g693(.A1(new_n890_), .A2(new_n711_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT61), .B(G155gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n890_), .B2(new_n264_), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n440_), .B(new_n377_), .C1(new_n838_), .C2(new_n848_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n899_), .A2(new_n251_), .A3(new_n259_), .A4(new_n580_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(KEYINPUT123), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n898_), .A2(new_n903_), .A3(new_n900_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1347gat));
  XOR2_X1   g704(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n441_), .A2(new_n655_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n908_), .A2(new_n668_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n857_), .A2(new_n638_), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n907_), .B1(new_n910_), .B2(new_n630_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n308_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n857_), .A2(new_n909_), .ZN(new_n913_));
  OAI211_X1 g712(.A(G169gat), .B(new_n906_), .C1(new_n913_), .C2(new_n639_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n912_), .A3(new_n914_), .ZN(G1348gat));
  INV_X1    g714(.A(new_n913_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n523_), .B1(new_n916_), .B2(new_n622_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n571_), .B1(new_n838_), .B2(new_n848_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n918_), .A2(G176gat), .A3(new_n622_), .A4(new_n908_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT125), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n920_), .ZN(G1349gat));
  AOI21_X1  g720(.A(new_n799_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n918_), .A2(new_n295_), .A3(new_n908_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n318_), .A2(new_n319_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n916_), .A2(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n913_), .B2(new_n264_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n259_), .A2(new_n327_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n913_), .B2(new_n927_), .ZN(G1351gat));
  XNOR2_X1  g727(.A(KEYINPUT127), .B(G197gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n655_), .A2(new_n577_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n859_), .A2(new_n662_), .A3(new_n571_), .A4(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n889_), .A2(KEYINPUT126), .A3(new_n571_), .A4(new_n930_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n929_), .B1(new_n935_), .B2(new_n638_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n929_), .ZN(new_n937_));
  AOI211_X1 g736(.A(new_n639_), .B(new_n937_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1352gat));
  AOI21_X1  g738(.A(G204gat), .B1(new_n935_), .B2(new_n622_), .ZN(new_n940_));
  AOI211_X1 g739(.A(new_n448_), .B(new_n740_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1353gat));
  OR2_X1    g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(new_n935_), .B2(new_n294_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT63), .B(G211gat), .ZN(new_n945_));
  AOI211_X1 g744(.A(new_n799_), .B(new_n945_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1354gat));
  AOI21_X1  g746(.A(G218gat), .B1(new_n935_), .B2(new_n259_), .ZN(new_n948_));
  INV_X1    g747(.A(G218gat), .ZN(new_n949_));
  AOI211_X1 g748(.A(new_n949_), .B(new_n264_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1355gat));
endmodule


