//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n208_), .B(new_n211_), .Z(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G229gat), .A3(G233gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n208_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n208_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(new_n211_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G229gat), .A2(G233gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT80), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G113gat), .B(G141gat), .Z(new_n222_));
  XNOR2_X1  g021(.A(G169gat), .B(G197gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  INV_X1    g026(.A(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(G190gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n230_), .B(new_n231_), .C1(G183gat), .C2(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G169gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(KEYINPUT86), .ZN(new_n239_));
  INV_X1    g038(.A(G176gat), .ZN(new_n240_));
  INV_X1    g039(.A(G169gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n241_), .A2(KEYINPUT22), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n240_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n232_), .B(new_n237_), .C1(new_n239_), .C2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n230_), .A2(new_n231_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n240_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT24), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n235_), .A2(new_n247_), .A3(KEYINPUT24), .A4(new_n236_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT84), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n254_), .A2(KEYINPUT84), .A3(new_n235_), .A4(new_n236_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT25), .B1(new_n228_), .B2(KEYINPUT81), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(G183gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n229_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n256_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT82), .B1(new_n229_), .B2(KEYINPUT26), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT26), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(G190gat), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n252_), .A2(new_n255_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n249_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(new_n255_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n264_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n268_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n245_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G99gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n271_), .B(KEYINPUT30), .ZN(new_n275_));
  INV_X1    g074(.A(G99gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G15gat), .B(G43gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT87), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(G71gat), .Z(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n274_), .A2(new_n277_), .A3(new_n285_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT90), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G134gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G127gat), .ZN(new_n291_));
  INV_X1    g090(.A(G127gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G134gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G120gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G113gat), .ZN(new_n296_));
  INV_X1    g095(.A(G113gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G120gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n291_), .A2(new_n293_), .A3(new_n296_), .A4(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n302_), .B(KEYINPUT31), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n289_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n287_), .A2(KEYINPUT90), .A3(new_n288_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n303_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(KEYINPUT1), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT91), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(G155gat), .A4(G162gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT91), .B1(new_n311_), .B2(KEYINPUT1), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G141gat), .B(G148gat), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT92), .A2(KEYINPUT3), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI22_X1  g122(.A1(KEYINPUT92), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n323_), .A2(new_n324_), .A3(new_n327_), .A4(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G155gat), .B(G162gat), .Z(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n320_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n302_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n318_), .A2(new_n319_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n302_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n336_), .A3(KEYINPUT4), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n302_), .B1(new_n320_), .B2(new_n331_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT100), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT100), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n337_), .A2(new_n344_), .A3(new_n338_), .A4(new_n341_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G85gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(KEYINPUT0), .B(G57gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n338_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n334_), .A2(new_n336_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n352_), .A3(KEYINPUT99), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT99), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n320_), .A2(new_n331_), .A3(new_n302_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n355_), .A2(new_n339_), .A3(new_n338_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n356_), .B2(new_n349_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n343_), .A2(new_n345_), .A3(new_n353_), .A4(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n338_), .B1(new_n355_), .B2(new_n339_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n335_), .A2(KEYINPUT4), .A3(new_n302_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n355_), .A2(new_n339_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(KEYINPUT4), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(new_n338_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n359_), .B1(new_n364_), .B2(new_n349_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n338_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n360_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n359_), .B(new_n349_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n358_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G8gat), .B(G36gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT18), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G197gat), .A2(G204gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT21), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383_));
  INV_X1    g182(.A(KEYINPUT94), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT21), .A3(new_n378_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT94), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n381_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(G190gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n254_), .A2(new_n233_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n246_), .A2(new_n396_), .A3(new_n248_), .A4(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n238_), .A2(new_n240_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n232_), .A2(new_n237_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n393_), .B2(new_n401_), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n377_), .B(new_n402_), .C1(new_n271_), .C2(new_n393_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n377_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n382_), .A2(new_n383_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n389_), .A2(new_n385_), .B1(new_n405_), .B2(new_n391_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n245_), .B(new_n406_), .C1(new_n267_), .C2(new_n270_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT20), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n393_), .B2(new_n401_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n404_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n375_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n271_), .A2(new_n393_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n402_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n404_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n377_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n416_), .A3(new_n374_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT101), .B1(new_n370_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n349_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT33), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n357_), .A2(new_n345_), .A3(new_n353_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n421_), .A2(new_n368_), .B1(new_n422_), .B2(new_n343_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT101), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n417_), .A4(new_n411_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n374_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n414_), .A2(new_n416_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT102), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n364_), .B(new_n349_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n414_), .A2(new_n416_), .A3(KEYINPUT102), .A4(new_n426_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n407_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n402_), .B1(new_n271_), .B2(new_n393_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n433_), .B2(new_n404_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT32), .A3(new_n374_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .A4(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n419_), .A2(new_n425_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n393_), .B(new_n438_), .C1(new_n439_), .C2(new_n335_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n438_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n320_), .B2(new_n331_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n406_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(KEYINPUT97), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT28), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n335_), .B2(new_n439_), .ZN(new_n448_));
  AND4_X1   g247(.A1(new_n447_), .A2(new_n320_), .A3(new_n331_), .A4(new_n439_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G22gat), .B(G50gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT28), .B1(new_n332_), .B2(KEYINPUT29), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n335_), .A2(new_n447_), .A3(new_n439_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n445_), .A2(KEYINPUT97), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n440_), .A2(new_n443_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n446_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n440_), .A2(new_n443_), .A3(KEYINPUT95), .A4(new_n445_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n451_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(new_n454_), .A3(new_n450_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n461_), .A2(KEYINPUT93), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT93), .B1(new_n461_), .B2(new_n462_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n440_), .A2(new_n443_), .A3(KEYINPUT95), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT95), .B1(new_n440_), .B2(new_n443_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n445_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n465_), .A2(new_n468_), .A3(KEYINPUT96), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n470_));
  AND4_X1   g269(.A1(KEYINPUT95), .A2(new_n440_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT93), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n467_), .A2(new_n445_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n440_), .A2(new_n443_), .A3(KEYINPUT95), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n470_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n459_), .B1(new_n469_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT98), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT96), .B1(new_n465_), .B2(new_n468_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n475_), .A2(new_n478_), .A3(new_n470_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT98), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(new_n459_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n437_), .A2(KEYINPUT103), .A3(new_n481_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT104), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n430_), .B(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n417_), .A2(KEYINPUT27), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n374_), .B(KEYINPUT105), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n434_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n490_), .A2(new_n492_), .B1(new_n418_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n485_), .B1(new_n484_), .B2(new_n459_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n459_), .ZN(new_n496_));
  AOI211_X1 g295(.A(KEYINPUT98), .B(new_n496_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n489_), .B(new_n494_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n487_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n495_), .A2(new_n497_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT103), .B1(new_n500_), .B2(new_n437_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n310_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n308_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n503_), .A2(new_n500_), .A3(new_n489_), .A4(new_n494_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n226_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G85gat), .ZN(new_n506_));
  INV_X1    g305(.A(G92gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT9), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G85gat), .B(G92gat), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n510_), .B2(KEYINPUT64), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT64), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n512_), .A3(KEYINPUT9), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT6), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n511_), .A2(new_n513_), .A3(new_n515_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n514_), .A2(KEYINPUT6), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n514_), .A2(KEYINPUT6), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(KEYINPUT66), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n276_), .A2(new_n517_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n522_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n520_), .B1(new_n529_), .B2(new_n509_), .ZN(new_n530_));
  AOI211_X1 g329(.A(KEYINPUT8), .B(new_n510_), .C1(new_n528_), .C2(new_n515_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n519_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT67), .B(G71gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G78gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n535_), .B(KEYINPUT11), .Z(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT68), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n532_), .A2(new_n539_), .A3(new_n543_), .A4(KEYINPUT12), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G230gat), .A2(G233gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT12), .B1(new_n532_), .B2(new_n539_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n540_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n532_), .A2(new_n539_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n550_), .B2(new_n540_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G120gat), .B(G148gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT5), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n549_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT70), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n542_), .A2(new_n544_), .B1(new_n540_), .B2(new_n547_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n551_), .B1(new_n559_), .B2(new_n546_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n556_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n560_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n556_), .B(KEYINPUT69), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT13), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n563_), .A2(KEYINPUT13), .A3(new_n566_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n208_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(new_n539_), .Z(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G155gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT17), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT79), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n574_), .A2(new_n582_), .A3(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n532_), .A2(new_n214_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n532_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT73), .A3(new_n211_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT73), .B1(new_n592_), .B2(new_n211_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n591_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n590_), .A2(new_n586_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n593_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n591_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G190gat), .B(G218gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT74), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT75), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n598_), .A2(new_n602_), .A3(KEYINPUT75), .A4(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n598_), .A2(new_n602_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n606_), .B(KEYINPUT36), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT76), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT37), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n608_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n505_), .A2(new_n571_), .A3(new_n585_), .A4(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT106), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n489_), .B(KEYINPUT107), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n203_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n618_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n569_), .A2(new_n570_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n631_), .A2(new_n226_), .A3(new_n584_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n489_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n626_), .A2(new_n627_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(new_n494_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n623_), .A2(new_n204_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT108), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n633_), .B2(new_n494_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n630_), .A2(KEYINPUT108), .A3(new_n637_), .A4(new_n632_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(G8gat), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT109), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(new_n644_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n638_), .B(new_n645_), .C1(new_n642_), .C2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n633_), .B2(new_n310_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT41), .Z(new_n651_));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n623_), .A2(new_n652_), .A3(new_n503_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  INV_X1    g454(.A(new_n500_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n623_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G22gat), .B1(new_n633_), .B2(new_n500_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1327gat));
  NAND2_X1  g459(.A1(new_n629_), .A2(new_n584_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT112), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(new_n571_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n505_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT113), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(KEYINPUT113), .A3(new_n505_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n489_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n571_), .A2(new_n225_), .A3(new_n584_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n571_), .A2(KEYINPUT110), .A3(new_n225_), .A4(new_n584_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n502_), .A2(new_n504_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n629_), .A2(new_n619_), .B1(new_n616_), .B2(KEYINPUT37), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT43), .B(new_n621_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n676_), .B(KEYINPUT44), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n625_), .A2(G29gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n671_), .B1(new_n687_), .B2(new_n688_), .ZN(G1328gat));
  NOR2_X1   g488(.A1(new_n494_), .A2(G36gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n666_), .A2(new_n667_), .A3(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n685_), .A2(new_n637_), .A3(new_n686_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT114), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(G36gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n693_), .B2(G36gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT46), .B(new_n692_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n687_), .A2(G43gat), .A3(new_n503_), .ZN(new_n702_));
  INV_X1    g501(.A(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n668_), .B2(new_n310_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g505(.A(G50gat), .B1(new_n669_), .B2(new_n656_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n656_), .A2(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n687_), .B2(new_n708_), .ZN(G1331gat));
  NOR2_X1   g508(.A1(new_n571_), .A2(new_n225_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n630_), .A2(new_n585_), .A3(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(new_n489_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n679_), .A2(new_n710_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n585_), .A3(new_n621_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n624_), .A2(G57gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n712_), .B1(new_n714_), .B2(new_n715_), .ZN(G1332gat));
  OAI21_X1  g515(.A(G64gat), .B1(new_n711_), .B2(new_n494_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n494_), .A2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n714_), .B2(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n711_), .B2(new_n310_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n310_), .A2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n714_), .B2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n711_), .B2(new_n500_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n500_), .A2(G78gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n714_), .B2(new_n728_), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n681_), .A2(new_n682_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT116), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n571_), .A2(new_n225_), .A3(new_n585_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT116), .B1(new_n681_), .B2(new_n682_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n489_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n713_), .A2(new_n662_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n506_), .A3(new_n625_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n737_), .B2(new_n637_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT117), .Z(new_n741_));
  NOR3_X1   g540(.A1(new_n735_), .A2(new_n507_), .A3(new_n494_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n735_), .B2(new_n310_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n503_), .A2(new_n516_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT118), .B1(new_n737_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g547(.A1(new_n733_), .A2(new_n656_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G106gat), .B1(new_n730_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT52), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n517_), .A3(new_n656_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(G1339gat));
  NAND4_X1  g554(.A1(new_n571_), .A2(new_n621_), .A3(new_n226_), .A4(new_n585_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n756_), .B(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n221_), .A2(new_n224_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n219_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n215_), .A2(new_n217_), .A3(new_n761_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n224_), .B(new_n762_), .C1(new_n212_), .C2(new_n219_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n563_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT121), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n549_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n559_), .A2(new_n546_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n768_), .B1(new_n549_), .B2(new_n767_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n565_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n549_), .A2(new_n767_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(new_n770_), .A3(new_n769_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n565_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n766_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n773_), .A2(new_n774_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n565_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n765_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n782_), .A2(new_n680_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n563_), .A2(new_n225_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n567_), .A2(new_n764_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n618_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT57), .B(new_n618_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n787_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n759_), .B1(new_n795_), .B2(new_n585_), .ZN(new_n796_));
  NOR4_X1   g595(.A1(new_n310_), .A2(new_n624_), .A3(new_n656_), .A4(new_n637_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT122), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n680_), .B1(new_n785_), .B2(KEYINPUT58), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n781_), .B(new_n765_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n782_), .A2(new_n786_), .A3(KEYINPUT122), .A4(new_n680_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n793_), .A4(new_n794_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n584_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n798_), .B1(new_n807_), .B2(new_n759_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n800_), .B(new_n225_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(G113gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(KEYINPUT123), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT123), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n756_), .B(new_n757_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n584_), .B2(new_n806_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n815_), .B2(new_n798_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n812_), .A2(new_n816_), .A3(new_n297_), .A4(new_n225_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n811_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT124), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n811_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1340gat));
  AND2_X1   g621(.A1(new_n812_), .A2(new_n816_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n295_), .B1(new_n571_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n823_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n295_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n800_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n826_));
  OAI21_X1  g625(.A(G120gat), .B1(new_n826_), .B2(new_n571_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1341gat));
  NAND3_X1  g627(.A1(new_n823_), .A2(new_n292_), .A3(new_n585_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G127gat), .B1(new_n826_), .B2(new_n584_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1342gat));
  NAND3_X1  g630(.A1(new_n823_), .A2(new_n290_), .A3(new_n629_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G134gat), .B1(new_n826_), .B2(new_n621_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1343gat));
  NAND2_X1  g633(.A1(new_n807_), .A2(new_n759_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n310_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n500_), .A2(new_n637_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n625_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n225_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n631_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n585_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  NOR2_X1   g645(.A1(new_n815_), .A2(new_n503_), .ZN(new_n847_));
  INV_X1    g646(.A(G162gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n838_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n629_), .A4(new_n849_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n836_), .A2(new_n621_), .A3(new_n838_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n848_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT125), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n850_), .B(KEYINPUT125), .C1(new_n851_), .C2(new_n848_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1347gat));
  NOR3_X1   g655(.A1(new_n625_), .A2(new_n310_), .A3(new_n494_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(new_n500_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n796_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n226_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT126), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT126), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n859_), .B2(new_n226_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(G169gat), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n861_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n860_), .A2(new_n238_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(G1348gat));
  NOR2_X1   g668(.A1(new_n815_), .A2(new_n656_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n857_), .A2(G176gat), .A3(new_n631_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n796_), .A2(new_n631_), .A3(new_n858_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n870_), .A2(new_n871_), .B1(new_n872_), .B2(new_n240_), .ZN(G1349gat));
  NOR3_X1   g672(.A1(new_n859_), .A2(new_n395_), .A3(new_n584_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n870_), .A2(new_n585_), .A3(new_n857_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n228_), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n859_), .B2(new_n621_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n629_), .A2(new_n394_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n859_), .B2(new_n878_), .ZN(G1351gat));
  NOR3_X1   g678(.A1(new_n500_), .A2(new_n670_), .A3(new_n494_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n847_), .A2(new_n225_), .A3(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g681(.A1(new_n847_), .A2(new_n880_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n571_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1353gat));
  NAND3_X1  g685(.A1(new_n847_), .A2(new_n585_), .A3(new_n880_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AND2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n887_), .B2(new_n888_), .ZN(G1354gat));
  OAI21_X1  g690(.A(G218gat), .B1(new_n883_), .B2(new_n621_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n618_), .A2(G218gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n883_), .B2(new_n893_), .ZN(G1355gat));
endmodule


