//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n967_, new_n968_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT93), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n204_), .A2(KEYINPUT93), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n207_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(new_n205_), .A3(new_n202_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT31), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT90), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT89), .B1(new_n223_), .B2(KEYINPUT22), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n222_), .B(new_n224_), .C1(new_n225_), .C2(KEYINPUT89), .ZN(new_n226_));
  AND3_X1   g025(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(new_n214_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n218_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT88), .A2(G169gat), .A3(G176gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n221_), .A2(new_n226_), .A3(new_n230_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n223_), .A3(new_n222_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n215_), .A2(new_n219_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n223_), .A2(new_n222_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n233_), .A2(new_n240_), .A3(KEYINPUT24), .A4(new_n234_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G190gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n217_), .A2(KEYINPUT26), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT25), .B1(new_n216_), .B2(KEYINPUT86), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT86), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(G183gat), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n248_), .B(new_n251_), .C1(new_n244_), .C2(new_n243_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n239_), .B(new_n241_), .C1(new_n247_), .C2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n236_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT30), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(G15gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(G43gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G71gat), .B(G99gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n256_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n254_), .B(KEYINPUT30), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n262_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT92), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n213_), .B1(new_n270_), .B2(KEYINPUT94), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(KEYINPUT94), .B2(new_n270_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G225gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n275_));
  INV_X1    g074(.A(G141gat), .ZN(new_n276_));
  INV_X1    g075(.A(G148gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n278_), .A2(KEYINPUT3), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT97), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n284_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT96), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n276_), .A4(new_n277_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT96), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n281_), .A2(new_n286_), .A3(new_n289_), .A4(new_n291_), .ZN(new_n292_));
  OR3_X1    g091(.A1(KEYINPUT95), .A2(G155gat), .A3(G162gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT95), .B1(G155gat), .B2(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT98), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT98), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n293_), .A2(new_n298_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n295_), .B(KEYINPUT1), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n294_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n278_), .B(new_n280_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n211_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n300_), .A2(new_n210_), .A3(new_n208_), .A4(new_n303_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(KEYINPUT106), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT106), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n308_), .A3(new_n211_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n275_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(KEYINPUT4), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n274_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n273_), .A3(new_n309_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G85gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT0), .B(G57gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n312_), .A2(new_n313_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n270_), .A2(KEYINPUT94), .A3(new_n212_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n272_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT103), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n300_), .A2(new_n325_), .A3(new_n303_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT28), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT99), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n300_), .A2(new_n329_), .A3(new_n325_), .A4(new_n303_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n328_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G22gat), .B(G50gat), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT99), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n334_), .B1(new_n338_), .B2(new_n331_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n324_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n304_), .A2(KEYINPUT29), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT100), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT21), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n344_), .A2(KEYINPUT21), .A3(new_n345_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n349_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n325_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(KEYINPUT100), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n343_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT101), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n359_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT102), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n353_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT102), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n341_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n363_), .B1(new_n343_), .B2(new_n356_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n361_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n335_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n338_), .A2(new_n334_), .A3(new_n331_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT103), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n340_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT103), .B1(new_n374_), .B2(new_n375_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n372_), .A3(new_n369_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT27), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT19), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n246_), .A2(new_n243_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT104), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n250_), .A2(new_n216_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT104), .B1(new_n391_), .B2(new_n386_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n385_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n240_), .A2(KEYINPUT24), .A3(new_n231_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n228_), .A2(new_n394_), .A3(new_n238_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT105), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n389_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(KEYINPUT104), .A3(new_n386_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n384_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n228_), .A2(new_n394_), .A3(new_n238_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT105), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n225_), .A2(new_n222_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n220_), .A3(new_n235_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n354_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT20), .B1(new_n254_), .B2(new_n353_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n383_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n354_), .A3(new_n405_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n254_), .B2(new_n353_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n383_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G8gat), .B(G36gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n408_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n408_), .B2(new_n413_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n381_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n417_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n406_), .A2(new_n407_), .A3(new_n383_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n393_), .A2(new_n395_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n365_), .A2(new_n423_), .A3(new_n366_), .A4(new_n405_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n412_), .B1(new_n411_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n421_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n408_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(KEYINPUT27), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n420_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n380_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n323_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n408_), .A2(new_n413_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n421_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n427_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n312_), .A2(new_n313_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n317_), .A2(KEYINPUT33), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n307_), .A2(new_n309_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT4), .ZN(new_n440_));
  INV_X1    g239(.A(new_n311_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n273_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT108), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT108), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n440_), .A2(new_n444_), .A3(new_n273_), .A4(new_n441_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT107), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n273_), .B1(new_n439_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n307_), .A2(KEYINPUT107), .A3(new_n309_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n317_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n443_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n438_), .B(new_n450_), .C1(KEYINPUT33), .C2(new_n320_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT109), .B1(new_n433_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n452_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OR3_X1    g254(.A1(new_n433_), .A2(KEYINPUT109), .A3(new_n452_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n455_), .B(new_n456_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n380_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n436_), .A2(new_n317_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n312_), .A2(new_n313_), .A3(new_n318_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n420_), .A4(new_n428_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT110), .B1(new_n380_), .B2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n377_), .A2(new_n379_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT110), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n429_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n272_), .A2(new_n322_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n432_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G113gat), .B(G141gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G169gat), .B(G197gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT85), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT78), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT79), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G1gat), .B(G8gat), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n477_), .A2(new_n483_), .A3(new_n481_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G29gat), .B(G36gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT73), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT73), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n487_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(new_n492_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n493_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT15), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n485_), .A2(new_n486_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT84), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT84), .B1(new_n507_), .B2(new_n508_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n499_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n496_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n498_), .B1(new_n497_), .B2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n474_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n509_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n497_), .B(new_n498_), .C1(new_n517_), .C2(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n474_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n515_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n470_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G85gat), .B(G92gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT10), .B(G99gat), .Z(new_n529_));
  INV_X1    g328(.A(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G85gat), .ZN(new_n532_));
  INV_X1    g331(.A(G92gat), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT9), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT64), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n526_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT6), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(G99gat), .A3(G106gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n528_), .A2(new_n531_), .A3(new_n536_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n538_), .A2(new_n540_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547_));
  INV_X1    g346(.A(G99gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n530_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n545_), .A2(new_n546_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT8), .B1(new_n552_), .B2(new_n526_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n549_), .A2(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n541_), .ZN(new_n555_));
  OR2_X1    g354(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n556_));
  NAND2_X1  g355(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n555_), .A2(new_n527_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n543_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(G71gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT67), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT67), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(G71gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(G78gat), .ZN(new_n565_));
  INV_X1    g364(.A(G78gat), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(G64gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(G57gat), .ZN(new_n569_));
  INV_X1    g368(.A(G57gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G64gat), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n569_), .A2(new_n571_), .A3(KEYINPUT11), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT11), .B1(new_n569_), .B2(new_n571_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n565_), .B(new_n567_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n569_), .A2(new_n571_), .A3(KEYINPUT11), .ZN(new_n575_));
  INV_X1    g374(.A(new_n567_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n566_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n575_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT68), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT68), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n525_), .B1(new_n559_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n546_), .A2(new_n551_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n538_), .A2(new_n540_), .A3(new_n544_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n526_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT8), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n558_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n581_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n574_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n590_), .B(new_n542_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n541_), .A2(KEYINPUT66), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n587_), .A3(new_n554_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n589_), .B1(new_n595_), .B2(new_n527_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n527_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n541_), .B2(new_n554_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n542_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n579_), .A2(KEYINPUT12), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n584_), .A2(new_n585_), .A3(new_n593_), .A4(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n585_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n559_), .A2(new_n583_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n592_), .A2(new_n591_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n599_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT72), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT70), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n608_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT13), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n608_), .A2(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n608_), .A2(new_n615_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(KEYINPUT13), .A3(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT76), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT34), .Z(new_n629_));
  INV_X1    g428(.A(KEYINPUT35), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT75), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n559_), .B2(new_n496_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n507_), .A2(new_n599_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n629_), .A2(new_n630_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n633_), .B(new_n634_), .C1(KEYINPUT74), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n632_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(KEYINPUT74), .C1(new_n599_), .C2(new_n513_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n599_), .B2(new_n513_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n542_), .A2(new_n590_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n639_), .B(new_n635_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n637_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n637_), .B2(new_n642_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n627_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT37), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n637_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(KEYINPUT77), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n646_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(G231gat), .ZN(new_n651_));
  INV_X1    g450(.A(G233gat), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n485_), .A2(new_n486_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n574_), .B(new_n578_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n654_), .A3(new_n579_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT68), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(new_n659_), .A3(new_n581_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G127gat), .B(G155gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(G183gat), .B(G211gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT17), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT17), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n661_), .A2(new_n662_), .A3(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n668_), .B(KEYINPUT81), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(new_n660_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT82), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT82), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n671_), .A2(new_n676_), .A3(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n650_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT83), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n524_), .A2(new_n622_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n321_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n478_), .A3(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT38), .ZN(new_n684_));
  INV_X1    g483(.A(new_n678_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n622_), .B2(new_n522_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n618_), .A2(new_n621_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n688_), .A2(KEYINPUT111), .A3(new_n523_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n646_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(KEYINPUT112), .B(new_n627_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n470_), .A2(new_n691_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n467_), .A2(new_n463_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n464_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n469_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n323_), .A2(new_n431_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n693_), .A2(new_n694_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT113), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n685_), .B(new_n690_), .C1(new_n696_), .C2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G1gat), .B1(new_n704_), .B2(new_n321_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n684_), .A2(new_n705_), .ZN(G1324gat));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n696_), .A2(new_n703_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n690_), .A2(new_n685_), .A3(new_n429_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n707_), .B(G8gat), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n691_), .B1(new_n470_), .B2(new_n695_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n701_), .A2(KEYINPUT113), .A3(new_n702_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT114), .B1(new_n713_), .B2(new_n479_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n710_), .A2(new_n714_), .A3(KEYINPUT39), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT39), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT114), .B(new_n716_), .C1(new_n713_), .C2(new_n479_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n681_), .A2(new_n479_), .A3(new_n429_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n715_), .A2(KEYINPUT40), .A3(new_n717_), .A4(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1325gat));
  INV_X1    g522(.A(new_n469_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n681_), .A2(new_n258_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G15gat), .B1(new_n704_), .B2(new_n469_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n726_), .A2(new_n727_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1326gat));
  INV_X1    g529(.A(G22gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n681_), .A2(new_n731_), .A3(new_n464_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G22gat), .B1(new_n704_), .B2(new_n380_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT42), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT42), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n734_), .B2(new_n735_), .ZN(G1327gat));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n646_), .B(new_n649_), .Z(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n470_), .B2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n701_), .A2(KEYINPUT43), .A3(new_n650_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n678_), .A3(new_n690_), .A4(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n701_), .A2(new_n650_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n685_), .B1(new_n744_), .B2(new_n737_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n745_), .A2(KEYINPUT44), .A3(new_n690_), .A4(new_n740_), .ZN(new_n746_));
  AND4_X1   g545(.A1(G29gat), .A2(new_n743_), .A3(new_n682_), .A4(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n678_), .A2(new_n695_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(new_n688_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n524_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G29gat), .B1(new_n751_), .B2(new_n682_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n747_), .A2(new_n752_), .ZN(G1328gat));
  NAND3_X1  g552(.A1(new_n743_), .A2(new_n746_), .A3(new_n429_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G36gat), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n430_), .A2(G36gat), .ZN(new_n756_));
  OR3_X1    g555(.A1(new_n750_), .A2(KEYINPUT45), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT45), .B1(new_n750_), .B2(new_n756_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(KEYINPUT46), .A3(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1329gat));
  NAND4_X1  g563(.A1(new_n743_), .A2(new_n746_), .A3(G43gat), .A4(new_n724_), .ZN(new_n765_));
  INV_X1    g564(.A(G43gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n750_), .B2(new_n469_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g568(.A1(G50gat), .A2(new_n743_), .A3(new_n464_), .A4(new_n746_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G50gat), .B1(new_n751_), .B2(new_n464_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1331gat));
  NAND2_X1  g571(.A1(new_n680_), .A2(new_n688_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n523_), .B(new_n701_), .C1(new_n773_), .C2(KEYINPUT115), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(KEYINPUT115), .B2(new_n773_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n570_), .A3(new_n682_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n675_), .A2(new_n677_), .A3(new_n523_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n622_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n696_), .B2(new_n703_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT116), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n778_), .C1(new_n696_), .C2(new_n703_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n780_), .A2(new_n682_), .A3(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n776_), .B1(new_n783_), .B2(new_n570_), .ZN(G1332gat));
  NAND3_X1  g583(.A1(new_n775_), .A2(new_n568_), .A3(new_n429_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n429_), .A3(new_n782_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G64gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G64gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1333gat));
  NAND3_X1  g589(.A1(new_n775_), .A2(new_n560_), .A3(new_n724_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n780_), .A2(new_n724_), .A3(new_n782_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(G71gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G71gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(G1334gat));
  NAND3_X1  g595(.A1(new_n775_), .A2(new_n566_), .A3(new_n464_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n780_), .A2(new_n464_), .A3(new_n782_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G78gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G78gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n622_), .A2(new_n522_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n739_), .A2(new_n678_), .A3(new_n740_), .A4(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n321_), .ZN(new_n805_));
  NOR4_X1   g604(.A1(new_n470_), .A2(new_n522_), .A3(new_n622_), .A4(new_n748_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n532_), .A3(new_n682_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT117), .Z(G1336gat));
  OAI21_X1  g608(.A(G92gat), .B1(new_n804_), .B2(new_n430_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n533_), .A3(new_n429_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1337gat));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n529_), .A3(new_n724_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT118), .ZN(new_n814_));
  OAI21_X1  g613(.A(G99gat), .B1(new_n804_), .B2(new_n469_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1338gat));
  NAND3_X1  g620(.A1(new_n806_), .A2(new_n530_), .A3(new_n464_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n823_), .B(G106gat), .C1(new_n804_), .C2(new_n380_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n745_), .A2(new_n464_), .A3(new_n740_), .A4(new_n803_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n823_), .B1(new_n826_), .B2(G106gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n822_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT53), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(new_n822_), .C1(new_n825_), .C2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1339gat));
  INV_X1    g631(.A(G113gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n523_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n614_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n608_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n498_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n497_), .B(new_n837_), .C1(new_n517_), .C2(new_n510_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n497_), .A2(new_n514_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n498_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n473_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n473_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n836_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n593_), .A2(new_n601_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n525_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n605_), .B2(new_n599_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n603_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT120), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n602_), .A2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n593_), .A2(new_n601_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT55), .A3(new_n585_), .A4(new_n584_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n854_), .B(new_n603_), .C1(new_n845_), .C2(new_n847_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n849_), .A2(new_n851_), .A3(new_n853_), .A4(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n614_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(KEYINPUT56), .A3(new_n614_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n844_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT58), .B1(new_n861_), .B2(KEYINPUT121), .ZN(new_n862_));
  INV_X1    g661(.A(new_n844_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n856_), .A2(KEYINPUT56), .A3(new_n614_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n614_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n862_), .A2(new_n650_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n522_), .A2(new_n836_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n841_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n843_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n616_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n702_), .C1(new_n872_), .C2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n702_), .B1(new_n872_), .B2(new_n877_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n516_), .A2(new_n521_), .B1(new_n608_), .B2(new_n835_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n876_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n886_), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n702_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n870_), .A2(new_n880_), .A3(new_n883_), .A4(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n678_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n688_), .A2(new_n777_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n738_), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n650_), .A2(new_n688_), .A3(new_n777_), .A4(KEYINPUT54), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n889_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  AOI21_X1  g696(.A(KEYINPUT59), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n431_), .A2(new_n321_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n878_), .A2(new_n879_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n695_), .B1(new_n885_), .B2(new_n876_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT122), .B1(new_n901_), .B2(KEYINPUT57), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n866_), .A2(new_n867_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n738_), .B1(new_n904_), .B2(KEYINPUT58), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n905_), .A2(new_n869_), .B1(new_n882_), .B2(new_n881_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n685_), .B1(new_n903_), .B2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n724_), .B(new_n899_), .C1(new_n907_), .C2(new_n894_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n898_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n894_), .B1(new_n888_), .B2(new_n678_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n899_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n469_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n910_), .B2(KEYINPUT123), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n834_), .B1(new_n909_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  AOI21_X1  g716(.A(G113gat), .B1(new_n912_), .B2(new_n522_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n917_), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n834_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n897_), .B1(new_n907_), .B2(new_n894_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n908_), .A2(new_n913_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n912_), .A2(new_n914_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n921_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT124), .B1(new_n925_), .B2(new_n918_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n920_), .A2(new_n926_), .ZN(G1340gat));
  INV_X1    g726(.A(G120gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n912_), .B(new_n929_), .C1(KEYINPUT60), .C2(new_n928_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n622_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n928_), .ZN(G1341gat));
  INV_X1    g731(.A(G127gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n912_), .A2(new_n933_), .A3(new_n685_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n678_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n933_), .ZN(G1342gat));
  INV_X1    g735(.A(G134gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n912_), .A2(new_n937_), .A3(new_n695_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n738_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n937_), .ZN(G1343gat));
  NAND2_X1  g739(.A1(new_n469_), .A2(new_n464_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n941_), .A2(new_n321_), .A3(new_n429_), .ZN(new_n942_));
  XOR2_X1   g741(.A(new_n942_), .B(KEYINPUT125), .Z(new_n943_));
  NAND2_X1  g742(.A1(new_n896_), .A2(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n523_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n276_), .ZN(G1344gat));
  NOR2_X1   g745(.A1(new_n944_), .A2(new_n622_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n277_), .ZN(G1345gat));
  NOR2_X1   g747(.A1(new_n944_), .A2(new_n678_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT61), .B(G155gat), .Z(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1346gat));
  OAI21_X1  g750(.A(G162gat), .B1(new_n944_), .B2(new_n738_), .ZN(new_n952_));
  OR2_X1    g751(.A1(new_n702_), .A2(G162gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n944_), .B2(new_n953_), .ZN(G1347gat));
  NOR2_X1   g753(.A1(new_n910_), .A2(new_n469_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n321_), .A2(new_n429_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n464_), .A2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n955_), .A2(new_n957_), .ZN(new_n958_));
  OAI21_X1  g757(.A(G169gat), .B1(new_n958_), .B2(new_n523_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n960_), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n955_), .A2(new_n522_), .A3(new_n225_), .A4(new_n957_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n961_), .A2(new_n962_), .A3(new_n963_), .ZN(G1348gat));
  NOR2_X1   g763(.A1(new_n958_), .A2(new_n622_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(new_n222_), .ZN(G1349gat));
  NOR2_X1   g765(.A1(new_n958_), .A2(new_n678_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n967_), .B1(new_n392_), .B2(new_n390_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n968_), .B1(new_n216_), .B2(new_n967_), .ZN(G1350gat));
  OAI21_X1  g768(.A(G190gat), .B1(new_n958_), .B2(new_n738_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n695_), .A2(new_n385_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n958_), .B2(new_n971_), .ZN(G1351gat));
  NOR3_X1   g771(.A1(new_n910_), .A2(new_n941_), .A3(new_n956_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(new_n522_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n688_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n678_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n973_), .A2(new_n978_), .A3(new_n979_), .ZN(new_n980_));
  INV_X1    g779(.A(new_n980_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n978_), .B1(new_n973_), .B2(new_n979_), .ZN(new_n982_));
  OAI22_X1  g781(.A1(new_n981_), .A2(new_n982_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n983_));
  INV_X1    g782(.A(new_n982_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n984_), .A2(new_n985_), .A3(new_n980_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n983_), .A2(new_n986_), .ZN(G1354gat));
  INV_X1    g786(.A(G218gat), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n973_), .A2(new_n988_), .A3(new_n695_), .ZN(new_n989_));
  AND2_X1   g788(.A1(new_n973_), .A2(new_n650_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n990_), .B2(new_n988_), .ZN(new_n991_));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  OAI211_X1 g792(.A(KEYINPUT127), .B(new_n989_), .C1(new_n990_), .C2(new_n988_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n993_), .A2(new_n994_), .ZN(G1355gat));
endmodule


