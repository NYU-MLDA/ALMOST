//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G85gat), .B(G92gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n208_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT66), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n219_), .A2(new_n214_), .A3(new_n215_), .A4(KEYINPUT65), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n211_), .A2(new_n213_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n223_));
  OAI211_X1 g022(.A(KEYINPUT8), .B(new_n204_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n217_), .A2(new_n212_), .A3(new_n220_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n204_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT64), .B(G92gat), .Z(new_n228_));
  INV_X1    g027(.A(G85gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT9), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n209_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT10), .B(G99gat), .Z(new_n232_));
  AOI22_X1  g031(.A1(KEYINPUT9), .A2(new_n204_), .B1(new_n232_), .B2(new_n215_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n225_), .A2(new_n227_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(KEYINPUT11), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n238_), .A3(KEYINPUT11), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n236_), .B2(KEYINPUT11), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n237_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT68), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n235_), .A4(new_n239_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n224_), .A2(new_n234_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n224_), .B2(new_n234_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n203_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n224_), .A2(new_n234_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n247_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n224_), .A2(new_n234_), .A3(new_n247_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n203_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT70), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G120gat), .B(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G176gat), .B(G204gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n254_), .A2(new_n260_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n203_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n257_), .A2(KEYINPUT12), .A3(new_n258_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(new_n252_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n266_), .B1(new_n271_), .B2(new_n259_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n268_), .A2(new_n272_), .A3(KEYINPUT71), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT71), .B1(new_n268_), .B2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n202_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n267_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n271_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n268_), .A2(new_n272_), .A3(KEYINPUT71), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT13), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n275_), .A2(KEYINPUT72), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT72), .B1(new_n275_), .B2(new_n281_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT73), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT73), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G29gat), .B(G36gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT15), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n255_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n224_), .A2(new_n234_), .A3(KEYINPUT75), .A4(new_n292_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G232gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT35), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n294_), .A2(new_n295_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT76), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n298_), .A2(new_n299_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n224_), .A2(new_n234_), .A3(new_n292_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .A4(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(new_n294_), .A3(new_n295_), .A4(new_n300_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n302_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT76), .B1(new_n298_), .B2(new_n299_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G190gat), .B(G218gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT77), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G134gat), .B(G162gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT36), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT78), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n316_), .B(KEYINPUT36), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n307_), .A2(new_n311_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(KEYINPUT79), .A3(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(KEYINPUT79), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT37), .A3(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT80), .B(KEYINPUT37), .Z(new_n326_));
  NAND3_X1  g125(.A1(new_n320_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n325_), .A2(KEYINPUT81), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT81), .B1(new_n325_), .B2(new_n327_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G231gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT83), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n247_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT82), .B(G8gat), .Z(new_n335_));
  INV_X1    g134(.A(G1gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT14), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G15gat), .B(G22gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G8gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n334_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n344_));
  XOR2_X1   g143(.A(G127gat), .B(G155gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G183gat), .B(G211gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n343_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n344_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n342_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n331_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n289_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT25), .B(G183gat), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT86), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G190gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT86), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(G183gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT25), .B(G183gat), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n359_), .B(new_n362_), .C1(new_n364_), .C2(new_n360_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT87), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(KEYINPUT24), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(KEYINPUT24), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT23), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(G183gat), .A3(G190gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n377_), .A3(KEYINPUT88), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n379_), .A3(KEYINPUT23), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n363_), .A2(new_n366_), .A3(new_n373_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(KEYINPUT89), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n374_), .A2(new_n384_), .A3(KEYINPUT23), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n385_), .A3(new_n377_), .ZN(new_n386_));
  OR2_X1    g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n389_));
  NOR3_X1   g188(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n382_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT30), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n382_), .A2(KEYINPUT30), .A3(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G43gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT90), .B(G15gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n399_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n397_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT91), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n397_), .A2(new_n398_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n407_), .B1(new_n406_), .B2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G127gat), .B(G134gat), .Z(new_n413_));
  XOR2_X1   g212(.A(G113gat), .B(G120gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT31), .Z(new_n416_));
  NOR2_X1   g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  AOI211_X1 g217(.A(new_n418_), .B(new_n407_), .C1(new_n406_), .C2(new_n411_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT105), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT103), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(KEYINPUT33), .ZN(new_n424_));
  INV_X1    g223(.A(new_n415_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  OR2_X1    g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT92), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT92), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(G141gat), .A3(G148gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT2), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(KEYINPUT95), .A2(KEYINPUT3), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n439_));
  OAI22_X1  g238(.A1(KEYINPUT95), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n426_), .B(new_n429_), .C1(new_n435_), .C2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n444_), .A2(new_n438_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n426_), .B1(new_n445_), .B2(new_n429_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n431_), .A2(new_n433_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n436_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n428_), .A2(KEYINPUT1), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT94), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n428_), .A2(new_n454_), .A3(KEYINPUT1), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n452_), .A2(new_n453_), .A3(new_n427_), .A4(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n428_), .A2(KEYINPUT1), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n427_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n454_), .B1(new_n428_), .B2(KEYINPUT1), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT94), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n450_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n425_), .B1(new_n447_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n429_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT96), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n457_), .A3(new_n456_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n450_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n465_), .A2(new_n442_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n415_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n469_), .A3(KEYINPUT4), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n442_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n466_), .A2(new_n467_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n415_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n471_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n472_), .A2(new_n473_), .A3(new_n415_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(new_n474_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n470_), .A2(new_n476_), .B1(new_n478_), .B2(new_n471_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G29gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G85gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n424_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n463_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n470_), .A2(new_n476_), .ZN(new_n487_));
  AND4_X1   g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n484_), .A4(new_n424_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G226gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n378_), .A2(new_n387_), .A3(new_n380_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT101), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n391_), .A2(new_n495_), .A3(new_n389_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n389_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT101), .B1(new_n497_), .B2(new_n390_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n500_));
  NOR2_X1   g299(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT100), .B(new_n372_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n368_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT100), .B1(new_n504_), .B2(new_n372_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n500_), .A2(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n367_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n364_), .A2(new_n359_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n386_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n499_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(G197gat), .A2(G204gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G197gat), .A2(G204gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(KEYINPUT21), .A3(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G211gat), .B(G218gat), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT21), .ZN(new_n518_));
  INV_X1    g317(.A(new_n514_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n512_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n515_), .A2(new_n520_), .A3(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT20), .B1(new_n511_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n382_), .B2(new_n392_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n493_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n382_), .A2(new_n524_), .A3(new_n392_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n511_), .A2(new_n522_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(KEYINPUT20), .A4(new_n492_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G8gat), .B(G36gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT18), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G64gat), .B(G92gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n530_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n471_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n463_), .A2(new_n469_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n484_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT104), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n470_), .B(new_n471_), .C1(KEYINPUT4), .C2(new_n463_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(KEYINPUT104), .A3(new_n538_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n535_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n422_), .B1(new_n489_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n487_), .A2(new_n486_), .A3(new_n484_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n424_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n479_), .A2(new_n484_), .A3(new_n424_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n551_), .A2(KEYINPUT105), .A3(new_n535_), .A4(new_n544_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n525_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n522_), .B1(new_n511_), .B2(KEYINPUT106), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n364_), .A2(new_n359_), .B1(new_n507_), .B2(new_n367_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n556_), .B(new_n386_), .C1(new_n505_), .C2(new_n503_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT106), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n499_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n554_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n553_), .B1(new_n560_), .B2(KEYINPUT107), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT107), .ZN(new_n562_));
  AOI211_X1 g361(.A(new_n562_), .B(new_n554_), .C1(new_n555_), .C2(new_n559_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n492_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n527_), .A2(new_n528_), .A3(KEYINPUT20), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(new_n492_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n534_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT32), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT108), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n547_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n487_), .A2(new_n486_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n538_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n487_), .A2(KEYINPUT108), .A3(new_n486_), .A4(new_n484_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n530_), .A2(new_n570_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n546_), .A2(new_n552_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT29), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n468_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT28), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(KEYINPUT28), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G228gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT97), .Z(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n585_), .A2(new_n586_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G22gat), .B(G50gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n522_), .B1(new_n468_), .B2(new_n582_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(G78gat), .ZN(new_n596_));
  INV_X1    g395(.A(G78gat), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n597_), .B(new_n522_), .C1(new_n468_), .C2(new_n582_), .ZN(new_n598_));
  AOI21_X1  g397(.A(G106gat), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(G106gat), .A3(new_n598_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n594_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n603_), .A2(new_n599_), .A3(new_n593_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n592_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n593_), .B1(new_n603_), .B2(new_n599_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n590_), .A2(new_n591_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n600_), .A2(new_n601_), .A3(new_n594_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n581_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n535_), .A2(KEYINPUT27), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT109), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n569_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n530_), .A2(new_n569_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT27), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n614_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n557_), .A2(new_n558_), .A3(new_n499_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n558_), .B1(new_n557_), .B2(new_n499_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n522_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n562_), .B1(new_n622_), .B2(new_n554_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n560_), .A2(KEYINPUT107), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n553_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n566_), .B1(new_n625_), .B2(new_n492_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT109), .B(new_n619_), .C1(new_n626_), .C2(new_n569_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n613_), .B1(new_n618_), .B2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n578_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n421_), .B1(new_n612_), .B2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n420_), .A2(new_n578_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n632_), .A2(new_n628_), .A3(new_n611_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n341_), .B(new_n292_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n341_), .A2(new_n293_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n636_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n341_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n292_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n637_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G113gat), .B(G141gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G169gat), .B(G197gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n643_), .B(new_n644_), .Z(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT85), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n642_), .B(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n634_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n578_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(G1gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n355_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT112), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n632_), .A2(new_n628_), .A3(new_n611_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n581_), .A2(new_n611_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(new_n421_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n320_), .A2(new_n322_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT111), .ZN(new_n662_));
  INV_X1    g461(.A(new_n353_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n661_), .B2(KEYINPUT111), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT72), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n273_), .A2(new_n274_), .A3(new_n202_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT13), .B1(new_n279_), .B2(new_n280_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n282_), .A3(new_n648_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT110), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n669_), .A2(new_n672_), .A3(new_n282_), .A4(new_n648_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n665_), .A2(new_n578_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G1gat), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n653_), .A2(new_n654_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n656_), .A2(new_n676_), .A3(new_n677_), .ZN(G1324gat));
  INV_X1    g477(.A(new_n628_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n662_), .A2(new_n664_), .A3(new_n674_), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT39), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(G8gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n680_), .B2(G8gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n355_), .A2(new_n650_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n679_), .A2(new_n335_), .ZN(new_n685_));
  OAI22_X1  g484(.A1(new_n682_), .A2(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1325gat));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n665_), .A2(new_n674_), .A3(new_n421_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(G15gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n690_), .B2(G15gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n689_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n694_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT41), .A3(new_n692_), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n684_), .A2(G15gat), .A3(new_n420_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n697_), .A3(new_n698_), .ZN(G1326gat));
  OR3_X1    g498(.A1(new_n684_), .A2(G22gat), .A3(new_n611_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n665_), .A2(new_n674_), .A3(new_n610_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G22gat), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT42), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT42), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1327gat));
  INV_X1    g504(.A(new_n285_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n353_), .A2(new_n660_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n650_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G29gat), .B1(new_n711_), .B2(new_n578_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n671_), .A2(new_n673_), .A3(new_n663_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n330_), .C1(new_n631_), .C2(new_n633_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n659_), .B2(new_n330_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n713_), .B(KEYINPUT44), .C1(new_n716_), .C2(new_n717_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n578_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n712_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  NOR2_X1   g523(.A1(KEYINPUT116), .A2(KEYINPUT46), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n628_), .A2(G36gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n728_));
  OR3_X1    g527(.A1(new_n710_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n710_), .B2(new_n727_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n720_), .A2(new_n679_), .A3(new_n721_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G36gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G36gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(KEYINPUT116), .A2(KEYINPUT46), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT117), .Z(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n731_), .B(new_n738_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1329gat));
  NAND3_X1  g541(.A1(new_n722_), .A2(G43gat), .A3(new_n421_), .ZN(new_n743_));
  INV_X1    g542(.A(G43gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n710_), .B2(new_n420_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g546(.A(G50gat), .B1(new_n711_), .B2(new_n610_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n610_), .A2(G50gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n722_), .B2(new_n749_), .ZN(G1331gat));
  NAND2_X1  g549(.A1(new_n659_), .A2(new_n649_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n751_), .A2(new_n354_), .A3(new_n285_), .ZN(new_n752_));
  INV_X1    g551(.A(G57gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n578_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n288_), .A2(new_n648_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n665_), .A2(new_n578_), .A3(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n756_), .B2(new_n753_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n758_), .A3(new_n679_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n755_), .A2(new_n662_), .A3(new_n679_), .A4(new_n664_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G64gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G64gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT118), .ZN(G1333gat));
  INV_X1    g564(.A(G71gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n752_), .A2(new_n766_), .A3(new_n421_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n665_), .A2(new_n421_), .A3(new_n755_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G71gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G71gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1334gat));
  NAND3_X1  g571(.A1(new_n752_), .A2(new_n597_), .A3(new_n610_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n665_), .A2(new_n610_), .A3(new_n755_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G78gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1335gat));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n634_), .B2(new_n331_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n715_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n648_), .A2(new_n353_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n706_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n651_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n288_), .A2(new_n708_), .A3(new_n751_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n229_), .A3(new_n578_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1336gat));
  AOI21_X1  g586(.A(G92gat), .B1(new_n785_), .B2(new_n679_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n679_), .A2(new_n228_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n782_), .B2(new_n789_), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n783_), .B2(new_n420_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n232_), .A3(new_n421_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g593(.A1(new_n782_), .A2(new_n610_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(G106gat), .A3(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n785_), .A2(new_n215_), .A3(new_n610_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n215_), .B1(new_n782_), .B2(new_n610_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT119), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n797_), .B(new_n798_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT53), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n799_), .A2(new_n801_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n797_), .A4(new_n798_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(G1339gat));
  AOI21_X1  g606(.A(new_n636_), .B1(new_n640_), .B2(new_n292_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n638_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n635_), .A2(new_n639_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n646_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n279_), .A2(new_n280_), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n270_), .A2(new_n269_), .A3(new_n252_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n254_), .A2(KEYINPUT55), .A3(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n266_), .C1(KEYINPUT55), .C2(new_n254_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n816_), .A2(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(KEYINPUT56), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n268_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n819_), .B2(new_n649_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n660_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n817_), .A2(new_n268_), .A3(new_n812_), .A4(new_n818_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n825_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n330_), .A3(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n820_), .B(new_n660_), .C1(KEYINPUT120), .C2(KEYINPUT57), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n823_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n648_), .B1(new_n275_), .B2(new_n281_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n353_), .B(new_n831_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n830_), .A2(new_n663_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n628_), .A2(new_n611_), .A3(new_n421_), .A4(new_n578_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n648_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n649_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n842_), .B2(new_n838_), .ZN(G1340gat));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n285_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n837_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n288_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n844_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n837_), .A2(new_n849_), .A3(new_n353_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n663_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n660_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n837_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n331_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n853_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n835_), .A2(new_n421_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n679_), .A2(new_n651_), .A3(new_n611_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n648_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n289_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g664(.A1(new_n860_), .A2(new_n663_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  OR3_X1    g667(.A1(new_n860_), .A2(G162gat), .A3(new_n660_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G162gat), .B1(new_n860_), .B2(new_n331_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1347gat));
  NOR2_X1   g670(.A1(new_n835_), .A2(new_n610_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n628_), .A2(new_n578_), .A3(new_n420_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n876_));
  AND2_X1   g675(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n875_), .B(new_n648_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n873_), .A2(new_n648_), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT121), .Z(new_n881_));
  NAND3_X1  g680(.A1(new_n872_), .A2(KEYINPUT122), .A3(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT122), .B1(new_n872_), .B2(new_n881_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n879_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(G169gat), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(new_n884_), .A3(KEYINPUT62), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n878_), .B1(new_n886_), .B2(new_n888_), .ZN(G1348gat));
  NAND3_X1  g688(.A1(new_n872_), .A2(new_n706_), .A3(new_n873_), .ZN(new_n890_));
  INV_X1    g689(.A(G176gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(KEYINPUT123), .A3(new_n891_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n872_), .A2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT124), .B1(new_n835_), .B2(new_n610_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n289_), .A2(G176gat), .A3(new_n873_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n894_), .A2(new_n895_), .B1(new_n899_), .B2(new_n900_), .ZN(G1349gat));
  NOR3_X1   g700(.A1(new_n874_), .A2(new_n364_), .A3(new_n663_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n873_), .A2(new_n353_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n897_), .A2(new_n903_), .A3(new_n898_), .A4(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(G183gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n897_), .A2(new_n898_), .A3(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT125), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n902_), .B1(new_n907_), .B2(new_n909_), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n874_), .B2(new_n331_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n854_), .A2(new_n359_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n874_), .B2(new_n912_), .ZN(G1351gat));
  NOR3_X1   g712(.A1(new_n611_), .A2(new_n628_), .A3(new_n578_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n858_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n649_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT126), .B(G197gat), .Z(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1352gat));
  INV_X1    g717(.A(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n289_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g720(.A1(new_n915_), .A2(new_n663_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT63), .B(G211gat), .Z(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n924_), .ZN(G1354gat));
  AOI21_X1  g724(.A(G218gat), .B1(new_n919_), .B2(new_n854_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n330_), .A2(G218gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT127), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n919_), .B2(new_n928_), .ZN(G1355gat));
endmodule


