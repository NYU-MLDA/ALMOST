//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  XNOR2_X1  g000(.A(KEYINPUT91), .B(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G228gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G155gat), .B(G162gat), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .A4(KEYINPUT89), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n205_), .B1(new_n214_), .B2(KEYINPUT89), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n204_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G155gat), .ZN(new_n217_));
  INV_X1    g016(.A(G162gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G155gat), .A3(G162gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n219_), .B(new_n221_), .C1(G155gat), .C2(G162gat), .ZN(new_n222_));
  XOR2_X1   g021(.A(G141gat), .B(G148gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n226_));
  INV_X1    g025(.A(G204gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G197gat), .ZN(new_n228_));
  INV_X1    g027(.A(G197gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G218gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G211gat), .ZN(new_n233_));
  INV_X1    g032(.A(G211gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G218gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n231_), .A2(new_n236_), .A3(KEYINPUT21), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G197gat), .B(G204gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n228_), .A2(new_n230_), .A3(new_n240_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n237_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n203_), .B1(new_n226_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n203_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n226_), .B2(KEYINPUT90), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n216_), .B2(new_n224_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT92), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n203_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n231_), .A2(KEYINPUT21), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n239_), .A2(new_n240_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n238_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n256_), .B2(new_n237_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT89), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT3), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n260_), .A2(new_n208_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n261_), .A2(new_n204_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n262_), .A2(KEYINPUT90), .A3(new_n248_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT92), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n258_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n245_), .B1(new_n252_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT90), .B1(new_n262_), .B2(new_n248_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n251_), .A2(new_n270_), .A3(KEYINPUT92), .A4(new_n257_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n267_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n245_), .A3(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G78gat), .B(G106gat), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n272_), .B2(new_n245_), .ZN(new_n278_));
  AOI211_X1 g077(.A(new_n244_), .B(new_n267_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n275_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G22gat), .B(G50gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT28), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n277_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G120gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G113gat), .ZN(new_n285_));
  INV_X1    g084(.A(G113gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G120gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G134gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G127gat), .ZN(new_n290_));
  INV_X1    g089(.A(G127gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G134gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n285_), .A2(new_n287_), .A3(new_n290_), .A4(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n225_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(KEYINPUT93), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT93), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n294_), .A2(new_n301_), .A3(new_n295_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n298_), .A2(new_n299_), .B1(new_n303_), .B2(new_n262_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n303_), .A2(new_n299_), .A3(new_n262_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n304_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT4), .B1(new_n304_), .B2(new_n305_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n296_), .B1(new_n216_), .B2(new_n224_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(KEYINPUT4), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n308_), .B1(new_n313_), .B2(new_n307_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G29gat), .ZN(new_n315_));
  INV_X1    g114(.A(G85gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT0), .B(G57gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n314_), .B(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n282_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n283_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n325_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT84), .B1(new_n325_), .B2(KEYINPUT23), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n324_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT83), .A3(G190gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n337_));
  INV_X1    g136(.A(G190gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT26), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n328_), .A2(new_n333_), .A3(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n325_), .A2(KEYINPUT23), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT86), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n325_), .A2(new_n345_), .A3(KEYINPUT23), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n342_), .B1(new_n347_), .B2(new_n324_), .ZN(new_n348_));
  INV_X1    g147(.A(G176gat), .ZN(new_n349_));
  AND2_X1   g148(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT85), .B(new_n349_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n332_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n341_), .B1(new_n348_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(G15gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n359_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n296_), .B(KEYINPUT31), .Z(new_n370_));
  OR2_X1    g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n367_), .A2(new_n368_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G92gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT18), .B(G64gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n357_), .A2(new_n243_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n243_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n346_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n345_), .B1(new_n325_), .B2(KEYINPUT23), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n324_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n389_));
  AND2_X1   g188(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n388_), .A2(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(new_n333_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n332_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT22), .B(G169gat), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n349_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n324_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n343_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n325_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n396_), .B1(new_n401_), .B2(new_n342_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n384_), .A2(new_n393_), .A3(new_n402_), .ZN(new_n403_));
  AND4_X1   g202(.A1(KEYINPUT20), .A2(new_n380_), .A3(new_n383_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n393_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(new_n243_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n394_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n397_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n355_), .B(new_n408_), .C1(new_n409_), .C2(new_n342_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n384_), .A2(new_n410_), .A3(new_n341_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n383_), .B1(new_n407_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n379_), .B1(new_n404_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n329_), .ZN(new_n414_));
  INV_X1    g213(.A(G169gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n349_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(KEYINPUT24), .A3(new_n332_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n392_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n409_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n352_), .A2(new_n332_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n342_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n328_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n243_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n411_), .A2(new_n423_), .A3(KEYINPUT20), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n382_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n379_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n380_), .A2(KEYINPUT20), .A3(new_n403_), .A4(new_n383_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n413_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT98), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT98), .ZN(new_n432_));
  AOI211_X1 g231(.A(new_n432_), .B(KEYINPUT27), .C1(new_n413_), .C2(new_n428_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(KEYINPUT27), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n380_), .A2(KEYINPUT20), .A3(new_n403_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n382_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n407_), .A2(new_n383_), .A3(new_n411_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n426_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT97), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n438_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n405_), .B1(new_n357_), .B2(new_n243_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n383_), .B1(new_n442_), .B2(new_n403_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n379_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(KEYINPUT27), .A4(new_n428_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n375_), .B1(new_n434_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n446_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n449_), .B(KEYINPUT99), .C1(new_n431_), .C2(new_n433_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n322_), .A2(new_n374_), .A3(new_n448_), .A4(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n282_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n276_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n278_), .A2(new_n279_), .A3(new_n275_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n277_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n320_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n431_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n429_), .A2(KEYINPUT98), .A3(new_n430_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n458_), .A2(new_n459_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT96), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n302_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n301_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI22_X1  g264(.A1(new_n465_), .A2(new_n225_), .B1(new_n310_), .B2(KEYINPUT94), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n303_), .A2(new_n299_), .A3(new_n262_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(KEYINPUT96), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n319_), .B1(new_n469_), .B2(new_n307_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n313_), .A2(new_n306_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n429_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n314_), .A2(new_n473_), .A3(KEYINPUT33), .A4(new_n319_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n307_), .B1(new_n476_), .B2(new_n311_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n308_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(KEYINPUT33), .A4(new_n319_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT95), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n319_), .A3(new_n478_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n472_), .A2(new_n474_), .A3(new_n480_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n425_), .A2(new_n485_), .A3(new_n427_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n441_), .A2(new_n443_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n487_), .A2(new_n485_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n314_), .A2(new_n319_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n481_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n486_), .B(new_n488_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n283_), .A2(new_n321_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n457_), .A2(new_n460_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n451_), .B1(new_n494_), .B2(new_n374_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G43gat), .B(G50gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(G29gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT82), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500_));
  INV_X1    g299(.A(G1gat), .ZN(new_n501_));
  INV_X1    g300(.A(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G1gat), .B(G8gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n499_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT81), .B(KEYINPUT15), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n498_), .B(new_n509_), .Z(new_n510_));
  MUX2_X1   g309(.A(new_n499_), .B(new_n510_), .S(new_n507_), .Z(new_n511_));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512_));
  MUX2_X1   g311(.A(new_n508_), .B(new_n511_), .S(new_n512_), .Z(new_n513_));
  XNOR2_X1  g312(.A(G113gat), .B(G141gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n513_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n495_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT100), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G85gat), .B(G92gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT6), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n526_), .B(new_n527_), .C1(G99gat), .C2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(G99gat), .ZN(new_n529_));
  INV_X1    g328(.A(G106gat), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n529_), .B(new_n530_), .C1(KEYINPUT68), .C2(KEYINPUT7), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT8), .B1(new_n523_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n525_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n532_), .B(KEYINPUT71), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n523_), .A2(KEYINPUT8), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n534_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n525_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT10), .B(G99gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT65), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n543_), .B2(new_n530_), .ZN(new_n544_));
  INV_X1    g343(.A(G92gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n316_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(KEYINPUT66), .A3(KEYINPUT9), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n316_), .A2(new_n545_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n547_), .B(new_n548_), .C1(new_n546_), .C2(KEYINPUT9), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT66), .B1(new_n546_), .B2(KEYINPUT9), .ZN(new_n550_));
  OR3_X1    g349(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT67), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT67), .B1(new_n549_), .B2(new_n550_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n544_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n540_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n510_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT79), .B(KEYINPUT34), .Z(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT35), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n555_), .B(new_n559_), .C1(new_n498_), .C2(new_n554_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(KEYINPUT35), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT80), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n560_), .A2(new_n563_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n564_), .A2(new_n565_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n568_), .B(KEYINPUT36), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n564_), .B2(new_n569_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT37), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n570_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT72), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n585_), .B2(KEYINPUT11), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n584_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT11), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n588_), .A2(new_n589_), .A3(new_n583_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n582_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n589_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n583_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n597_), .A3(new_n581_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n507_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n234_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT16), .B(G183gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT17), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(KEYINPUT17), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n604_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n580_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT78), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT64), .Z(new_n619_));
  NOR3_X1   g418(.A1(new_n591_), .A2(new_n582_), .A3(new_n592_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n581_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n540_), .A2(new_n553_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n554_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT12), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n593_), .A2(new_n598_), .B1(new_n553_), .B2(new_n540_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT12), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n593_), .A2(new_n598_), .A3(new_n553_), .A4(new_n540_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT75), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n623_), .A2(KEYINPUT75), .A3(new_n598_), .A4(new_n593_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n628_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n619_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n630_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(G176gat), .B(G204gat), .Z(new_n638_));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n637_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n630_), .B(new_n642_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(KEYINPUT77), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT77), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n637_), .A2(new_n647_), .A3(new_n643_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(KEYINPUT13), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT13), .B1(new_n646_), .B2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n617_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n648_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT13), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(KEYINPUT13), .A3(new_n648_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(KEYINPUT78), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n651_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n520_), .A2(new_n616_), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n501_), .A3(new_n320_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n661_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n492_), .A2(new_n493_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n455_), .A2(new_n456_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n320_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n460_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n374_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n448_), .A2(new_n374_), .A3(new_n450_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n493_), .A2(new_n666_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n571_), .A2(new_n574_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n672_), .A2(new_n615_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n654_), .A2(new_n655_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(KEYINPUT102), .A3(new_n518_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n649_), .A2(new_n650_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n518_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n676_), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G1gat), .B1(new_n681_), .B2(new_n666_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n662_), .A2(new_n663_), .A3(new_n682_), .ZN(G1324gat));
  NAND2_X1  g482(.A1(new_n448_), .A2(new_n450_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n659_), .A2(new_n502_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G8gat), .B1(new_n681_), .B2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(KEYINPUT103), .A3(KEYINPUT39), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(KEYINPUT39), .B2(new_n687_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT103), .B1(new_n687_), .B2(KEYINPUT39), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(G1325gat));
  INV_X1    g492(.A(new_n374_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G15gat), .B1(new_n681_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT41), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n659_), .A2(new_n361_), .A3(new_n374_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n681_), .B2(new_n493_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n659_), .A2(new_n701_), .A3(new_n665_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1327gat));
  INV_X1    g502(.A(G29gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n580_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n706_), .A3(KEYINPUT43), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n680_), .A2(new_n676_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n615_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n711_), .A2(new_n712_), .A3(KEYINPUT44), .A4(new_n615_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n320_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n704_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n718_), .B2(new_n717_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n615_), .A2(KEYINPUT106), .A3(new_n673_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722_));
  INV_X1    g521(.A(new_n673_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n614_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n678_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n520_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n320_), .A2(new_n704_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT107), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n720_), .B1(new_n728_), .B2(new_n730_), .ZN(G1328gat));
  NAND2_X1  g530(.A1(new_n715_), .A2(new_n716_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G36gat), .B1(new_n732_), .B2(new_n686_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n686_), .A2(G36gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n520_), .A2(new_n727_), .A3(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT45), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(KEYINPUT46), .A3(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1329gat));
  OAI21_X1  g540(.A(new_n363_), .B1(new_n728_), .B2(new_n694_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n374_), .A2(G43gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n732_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g544(.A(G50gat), .B1(new_n732_), .B2(new_n493_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n493_), .A2(G50gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT108), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n728_), .B2(new_n748_), .ZN(G1331gat));
  AND4_X1   g548(.A1(new_n679_), .A2(new_n616_), .A3(new_n495_), .A4(new_n678_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n320_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n518_), .B1(new_n651_), .B2(new_n656_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n674_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n320_), .A2(G57gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1332gat));
  INV_X1    g555(.A(G64gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n750_), .A2(new_n757_), .A3(new_n684_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G64gat), .B1(new_n753_), .B2(new_n686_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n761_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n758_), .B1(new_n762_), .B2(new_n763_), .ZN(G1333gat));
  INV_X1    g563(.A(G71gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n750_), .A2(new_n765_), .A3(new_n374_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G71gat), .B1(new_n753_), .B2(new_n694_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT49), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT49), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT110), .ZN(G1334gat));
  OAI21_X1  g570(.A(G78gat), .B1(new_n753_), .B2(new_n493_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT50), .ZN(new_n773_));
  INV_X1    g572(.A(G78gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n750_), .A2(new_n774_), .A3(new_n665_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1335gat));
  NOR3_X1   g575(.A1(new_n675_), .A2(new_n518_), .A3(new_n614_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n711_), .A2(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n778_), .A2(new_n316_), .A3(new_n666_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n726_), .A2(new_n672_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n752_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n320_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n779_), .A2(new_n782_), .ZN(G1336gat));
  OAI21_X1  g582(.A(G92gat), .B1(new_n778_), .B2(new_n686_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n545_), .A3(new_n684_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT111), .ZN(G1337gat));
  AND2_X1   g586(.A1(new_n374_), .A2(new_n543_), .ZN(new_n788_));
  AND4_X1   g587(.A1(new_n495_), .A2(new_n752_), .A3(new_n725_), .A4(new_n788_), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT104), .B(new_n708_), .C1(new_n495_), .C2(new_n580_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT43), .B1(new_n705_), .B2(new_n706_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n374_), .B(new_n777_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n792_), .B2(G99gat), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT113), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(G99gat), .ZN(new_n796_));
  INV_X1    g595(.A(new_n789_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n794_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n799_), .B(new_n789_), .C1(new_n792_), .C2(G99gat), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n795_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT51), .B1(new_n793_), .B2(KEYINPUT112), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n804_), .A2(new_n801_), .A3(KEYINPUT113), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT114), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n795_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n800_), .A2(new_n802_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n806_), .A2(new_n812_), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n781_), .A2(new_n530_), .A3(new_n665_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n711_), .A2(new_n665_), .A3(new_n777_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(G106gat), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n815_), .B2(G106gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g619(.A1(new_n518_), .A2(new_n645_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT75), .B1(new_n622_), .B2(new_n623_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n631_), .A2(new_n632_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n627_), .B(new_n629_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n619_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n624_), .A2(new_n627_), .A3(new_n629_), .A4(KEYINPUT55), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n630_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .A4(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n643_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n825_), .A2(new_n619_), .B1(new_n630_), .B2(new_n829_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n828_), .B1(new_n833_), .B2(new_n827_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n822_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n826_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT117), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n837_), .A2(KEYINPUT56), .A3(new_n643_), .A4(new_n831_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n821_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n513_), .A2(new_n517_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n512_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n508_), .A2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n842_), .B(new_n516_), .C1(new_n512_), .C2(new_n511_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT118), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n845_), .A2(new_n648_), .A3(new_n646_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n723_), .B1(new_n839_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT57), .B(new_n723_), .C1(new_n839_), .C2(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n845_), .A2(new_n645_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n853_), .A2(KEYINPUT58), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n580_), .B1(new_n853_), .B2(KEYINPUT58), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n615_), .B1(new_n851_), .B2(new_n856_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n579_), .A2(new_n679_), .A3(new_n614_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n675_), .A3(new_n859_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n860_), .A2(KEYINPUT116), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(KEYINPUT116), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n858_), .A2(new_n675_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n861_), .B(new_n862_), .C1(new_n859_), .C2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n666_), .B1(new_n857_), .B2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n669_), .A2(new_n665_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867_), .B2(new_n518_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n857_), .A2(new_n864_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n869_), .A2(KEYINPUT119), .A3(new_n320_), .A4(new_n866_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n865_), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n866_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n286_), .B1(new_n518_), .B2(KEYINPUT120), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(KEYINPUT120), .B2(new_n286_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n868_), .B1(new_n874_), .B2(new_n876_), .ZN(G1340gat));
  OAI21_X1  g676(.A(new_n284_), .B1(new_n675_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n867_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n284_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n658_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n284_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n867_), .B2(new_n614_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n615_), .A2(KEYINPUT121), .ZN(new_n883_));
  MUX2_X1   g682(.A(KEYINPUT121), .B(new_n883_), .S(G127gat), .Z(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n874_), .B2(new_n884_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n867_), .B2(new_n673_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n579_), .A2(new_n289_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n874_), .B2(new_n887_), .ZN(G1343gat));
  NAND3_X1  g687(.A1(new_n686_), .A2(new_n665_), .A3(new_n694_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n865_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n518_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT122), .B(G141gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n893_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n518_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n865_), .A2(new_n657_), .A3(new_n890_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT123), .B(G148gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n865_), .A2(new_n614_), .A3(new_n890_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  NAND3_X1  g702(.A1(new_n891_), .A2(G162gat), .A3(new_n580_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n865_), .A2(new_n673_), .A3(new_n890_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n906_), .A3(new_n218_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n905_), .B2(new_n218_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1347gat));
  XOR2_X1   g709(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n686_), .A2(new_n694_), .A3(new_n670_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n869_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n679_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n912_), .B1(new_n915_), .B2(new_n415_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n395_), .ZN(new_n917_));
  OAI211_X1 g716(.A(G169gat), .B(new_n911_), .C1(new_n914_), .C2(new_n679_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(G1348gat));
  NOR3_X1   g718(.A1(new_n914_), .A2(new_n349_), .A3(new_n658_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n914_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n678_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n349_), .B2(new_n922_), .ZN(G1349gat));
  NOR2_X1   g722(.A1(new_n914_), .A2(new_n615_), .ZN(new_n924_));
  MUX2_X1   g723(.A(G183gat), .B(new_n334_), .S(new_n924_), .Z(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n914_), .B2(new_n579_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n673_), .B1(new_n391_), .B2(new_n390_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n914_), .B2(new_n927_), .ZN(G1351gat));
  NAND2_X1  g727(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n684_), .A2(new_n457_), .A3(new_n694_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n869_), .A2(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n931_), .B2(new_n679_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n931_), .A2(new_n658_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n227_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AND2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  NOR4_X1   g737(.A1(new_n931_), .A2(new_n615_), .A3(new_n937_), .A4(new_n938_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n869_), .A2(new_n930_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n614_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n941_), .B2(new_n937_), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n940_), .B2(new_n673_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n580_), .A2(G218gat), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n931_), .A2(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(KEYINPUT127), .B1(new_n943_), .B2(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n232_), .B1(new_n931_), .B2(new_n723_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n947_), .B(new_n948_), .C1(new_n931_), .C2(new_n944_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n946_), .A2(new_n949_), .ZN(G1355gat));
endmodule


