//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n203_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT25), .B(G183gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(new_n212_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  OR3_X1    g016(.A1(new_n204_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT22), .B1(new_n204_), .B2(KEYINPUT81), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n205_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT82), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n214_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT30), .Z(new_n223_));
  NAND2_X1  g022(.A1(G227gat), .A2(G233gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT83), .ZN(new_n225_));
  XOR2_X1   g024(.A(G71gat), .B(G99gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G15gat), .B(G43gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n230_), .B(KEYINPUT84), .Z(new_n231_));
  NOR2_X1   g030(.A1(new_n223_), .A2(new_n229_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT85), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT87), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(G134gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT86), .B(G127gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(KEYINPUT31), .Z(new_n239_));
  OR2_X1    g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT22), .B(G169gat), .Z(new_n243_));
  OAI21_X1  g042(.A(new_n216_), .B1(G176gat), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT98), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n211_), .A2(new_n213_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT97), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n208_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n251_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT91), .ZN(new_n257_));
  INV_X1    g056(.A(new_n255_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT92), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT92), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n252_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n249_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT93), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n262_), .B(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n263_), .B(KEYINPUT20), .C1(new_n265_), .C2(new_n222_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n272_));
  INV_X1    g071(.A(new_n249_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n262_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n265_), .A2(new_n222_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n269_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G64gat), .B(G92gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT32), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT88), .Z(new_n289_));
  NAND2_X1  g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(G155gat), .B(G162gat), .Z(new_n291_));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n289_), .A2(new_n290_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT89), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n288_), .B(KEYINPUT3), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n290_), .B(KEYINPUT2), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT90), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n291_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(new_n238_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT4), .ZN(new_n305_));
  AOI211_X1 g104(.A(KEYINPUT4), .B(new_n238_), .C1(new_n297_), .C2(new_n302_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT100), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(KEYINPUT100), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n305_), .A2(new_n307_), .A3(new_n309_), .A4(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n304_), .A2(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G57gat), .B(G85gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G29gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n311_), .A2(new_n318_), .A3(new_n312_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n266_), .A2(new_n269_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n274_), .A2(new_n244_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n272_), .B1(new_n324_), .B2(new_n248_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n276_), .A3(new_n270_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n287_), .B(new_n322_), .C1(new_n286_), .C2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n321_), .B(KEYINPUT33), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n279_), .A2(new_n285_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n318_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT102), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n305_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n332_), .B1(new_n309_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n278_), .A2(new_n284_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n328_), .B1(new_n329_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n303_), .A2(KEYINPUT29), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n265_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT94), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n262_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT94), .B1(new_n303_), .B2(KEYINPUT29), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n340_), .B1(new_n344_), .B2(new_n338_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n346_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n303_), .A2(KEYINPUT29), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT28), .Z(new_n351_));
  XOR2_X1   g150(.A(G78gat), .B(G106gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT95), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n351_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n337_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n330_), .A2(new_n335_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n322_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n330_), .B(KEYINPUT27), .C1(new_n285_), .C2(new_n327_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n360_), .A2(new_n363_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n242_), .B1(new_n359_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n242_), .A2(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n365_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n360_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G29gat), .B(G36gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G43gat), .B(G50gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n374_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n372_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT15), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G15gat), .B(G22gat), .ZN(new_n381_));
  INV_X1    g180(.A(G1gat), .ZN(new_n382_));
  INV_X1    g181(.A(G8gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT14), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G1gat), .B(G8gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n380_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G229gat), .A2(G233gat), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n387_), .A2(new_n378_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n387_), .B(new_n378_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n389_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G113gat), .B(G141gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G169gat), .B(G197gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n391_), .A2(new_n394_), .A3(KEYINPUT79), .A4(new_n398_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n391_), .A2(new_n394_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n397_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(KEYINPUT80), .A3(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G230gat), .A2(G233gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT65), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(KEYINPUT65), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n413_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(KEYINPUT65), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(G99gat), .A4(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT66), .ZN(new_n422_));
  OAI22_X1  g221(.A1(new_n422_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT7), .ZN(new_n424_));
  INV_X1    g223(.A(G99gat), .ZN(new_n425_));
  INV_X1    g224(.A(G106gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .A4(KEYINPUT66), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n418_), .A2(new_n421_), .A3(new_n423_), .A4(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(G85gat), .A2(G92gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G85gat), .A2(G92gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(KEYINPUT68), .A3(new_n430_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n425_), .A2(KEYINPUT10), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G99gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT64), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n426_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n418_), .A2(new_n421_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n430_), .A2(KEYINPUT9), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n429_), .A2(KEYINPUT9), .A3(new_n430_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n449_), .A2(new_n450_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n438_), .A2(KEYINPUT67), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n440_), .A2(KEYINPUT67), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n428_), .A2(new_n435_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n441_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n460_));
  XOR2_X1   g259(.A(G71gat), .B(G78gat), .Z(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n459_), .B(KEYINPUT11), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n461_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(KEYINPUT70), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT70), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n441_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n464_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT71), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n470_), .A2(new_n471_), .B1(new_n468_), .B2(new_n467_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n465_), .A2(KEYINPUT71), .A3(new_n469_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n412_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT72), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n443_), .A2(G99gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n425_), .A2(KEYINPUT10), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT64), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(G106gat), .B1(new_n478_), .B2(new_n446_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n418_), .A2(new_n421_), .A3(new_n453_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n451_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n439_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n475_), .B1(new_n483_), .B2(new_n457_), .ZN(new_n484_));
  AND4_X1   g283(.A1(new_n475_), .A2(new_n441_), .A3(new_n454_), .A4(new_n457_), .ZN(new_n485_));
  OAI211_X1 g284(.A(KEYINPUT12), .B(new_n468_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n412_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n467_), .A2(new_n468_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT73), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT73), .ZN(new_n492_));
  AOI211_X1 g291(.A(new_n492_), .B(KEYINPUT12), .C1(new_n467_), .C2(new_n468_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n486_), .B(new_n488_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT5), .B(G176gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G204gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G120gat), .B(G148gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  OR3_X1    g298(.A1(new_n474_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(new_n474_), .B2(new_n495_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT74), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n503_), .B2(KEYINPUT13), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n371_), .A2(new_n411_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G190gat), .B(G218gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G134gat), .B(G162gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n467_), .B(KEYINPUT72), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT34), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n515_), .A2(new_n380_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n516_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n467_), .A2(new_n378_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT75), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n521_), .A2(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n520_), .A2(new_n529_), .A3(new_n523_), .A4(new_n525_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n514_), .B1(new_n531_), .B2(KEYINPUT76), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n533_), .B(new_n513_), .C1(new_n528_), .C2(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  OR3_X1    g335(.A1(new_n532_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT78), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(KEYINPUT37), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n532_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n540_), .B1(new_n541_), .B2(KEYINPUT78), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n387_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n464_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G127gat), .B(G155gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G211gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT16), .B(G183gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n549_), .A2(KEYINPUT17), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n549_), .A2(KEYINPUT17), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n545_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n539_), .A2(new_n542_), .A3(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n508_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n382_), .A3(new_n322_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT38), .ZN(new_n558_));
  INV_X1    g357(.A(new_n554_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n537_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n508_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(G1gat), .B1(new_n561_), .B2(new_n364_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(G1324gat));
  INV_X1    g362(.A(new_n369_), .ZN(new_n564_));
  OAI21_X1  g363(.A(G8gat), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n556_), .A2(new_n383_), .A3(new_n369_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT40), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(G1325gat));
  INV_X1    g370(.A(new_n242_), .ZN(new_n572_));
  OAI21_X1  g371(.A(G15gat), .B1(new_n561_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(G15gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n556_), .A2(new_n576_), .A3(new_n242_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT105), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(KEYINPUT105), .A3(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(G1326gat));
  OAI21_X1  g381(.A(G22gat), .B1(new_n561_), .B2(new_n358_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT42), .ZN(new_n584_));
  INV_X1    g383(.A(G22gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n556_), .A2(new_n585_), .A3(new_n360_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(G1327gat));
  NOR2_X1   g386(.A1(new_n507_), .A2(new_n411_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n541_), .A2(new_n554_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n588_), .B(new_n589_), .C1(new_n367_), .C2(new_n370_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(new_n364_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n539_), .A2(new_n542_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT43), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT43), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n559_), .B(new_n588_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT44), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n593_), .B(KEYINPUT43), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(KEYINPUT44), .A3(new_n559_), .A4(new_n588_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n322_), .A3(new_n600_), .ZN(new_n601_));
  MUX2_X1   g400(.A(new_n591_), .B(new_n601_), .S(G29gat), .Z(G1328gat));
  INV_X1    g401(.A(KEYINPUT46), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT107), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(KEYINPUT107), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n600_), .A3(new_n369_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G36gat), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n590_), .A2(G36gat), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT106), .B1(new_n608_), .B2(new_n564_), .ZN(new_n609_));
  OR4_X1    g408(.A1(KEYINPUT106), .A2(new_n590_), .A3(G36gat), .A4(new_n564_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n609_), .A2(new_n610_), .A3(KEYINPUT45), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT45), .B1(new_n609_), .B2(new_n610_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n604_), .B(new_n605_), .C1(new_n607_), .C2(new_n613_), .ZN(new_n614_));
  AND4_X1   g413(.A1(KEYINPUT107), .A2(new_n607_), .A3(new_n613_), .A4(new_n603_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1329gat));
  NAND4_X1  g415(.A1(new_n598_), .A2(new_n600_), .A3(G43gat), .A4(new_n242_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n590_), .A2(new_n572_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(G43gat), .B2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g419(.A1(new_n598_), .A2(new_n600_), .A3(G50gat), .A4(new_n360_), .ZN(new_n621_));
  INV_X1    g420(.A(G50gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n590_), .B2(new_n358_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1331gat));
  NAND2_X1  g423(.A1(new_n507_), .A2(new_n411_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n371_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n555_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G57gat), .B1(new_n627_), .B2(new_n322_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n560_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n364_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(G57gat), .B2(new_n630_), .ZN(G1332gat));
  OAI21_X1  g430(.A(G64gat), .B1(new_n629_), .B2(new_n564_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(G64gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n627_), .A2(new_n635_), .A3(new_n369_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(G1333gat));
  INV_X1    g436(.A(G71gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n627_), .A2(new_n638_), .A3(new_n242_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n629_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n640_), .B2(new_n242_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT49), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n642_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n639_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT109), .ZN(G1334gat));
  OAI21_X1  g446(.A(G78gat), .B1(new_n629_), .B2(new_n358_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT50), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n358_), .A2(G78gat), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT110), .Z(new_n651_));
  NAND2_X1  g450(.A1(new_n627_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(G1335gat));
  NAND2_X1  g452(.A1(new_n626_), .A2(new_n589_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G85gat), .B1(new_n655_), .B2(new_n322_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n625_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n599_), .A2(new_n559_), .A3(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n364_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n656_), .B1(new_n659_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g459(.A(G92gat), .B1(new_n655_), .B2(new_n369_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n658_), .A2(new_n564_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g462(.A(G99gat), .B1(new_n658_), .B2(new_n572_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n242_), .B1(new_n448_), .B2(new_n447_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n654_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g466(.A1(new_n655_), .A2(new_n426_), .A3(new_n360_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n599_), .A2(new_n559_), .A3(new_n360_), .A4(new_n657_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT52), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(G106gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G106gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g473(.A(KEYINPUT54), .ZN(new_n675_));
  INV_X1    g474(.A(new_n507_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n555_), .A2(new_n675_), .A3(new_n411_), .A4(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n539_), .A2(new_n542_), .A3(new_n554_), .A4(new_n411_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT54), .B1(new_n678_), .B2(new_n507_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT57), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n486_), .B(new_n470_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n487_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT55), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n494_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT12), .B1(new_n467_), .B2(new_n468_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT73), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n687_), .A2(KEYINPUT55), .A3(new_n488_), .A4(new_n486_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n685_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n499_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT112), .B(KEYINPUT56), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT113), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT56), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT114), .B1(new_n690_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT114), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n689_), .A2(new_n697_), .A3(KEYINPUT56), .A4(new_n499_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(KEYINPUT113), .A3(new_n691_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n694_), .A2(new_n696_), .A3(new_n698_), .A4(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT115), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n410_), .A2(new_n500_), .A3(KEYINPUT111), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT111), .B1(new_n410_), .B2(new_n500_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n700_), .A2(new_n701_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n701_), .B1(new_n700_), .B2(new_n704_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n388_), .A2(new_n393_), .A3(new_n390_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n392_), .A2(new_n389_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n397_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n403_), .A2(new_n709_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT116), .Z(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n502_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT117), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(KEYINPUT117), .A3(new_n502_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n705_), .A2(new_n706_), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n681_), .B1(new_n717_), .B2(new_n537_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n700_), .A2(new_n704_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT115), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n700_), .A2(new_n701_), .A3(new_n704_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT57), .B(new_n541_), .C1(new_n722_), .C2(new_n716_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n690_), .B(new_n695_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n500_), .A3(new_n711_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT58), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n592_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n718_), .A2(new_n723_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n680_), .B1(new_n728_), .B2(new_n559_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n369_), .A2(new_n360_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n572_), .A2(new_n364_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n729_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G113gat), .B1(new_n734_), .B2(new_n410_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT118), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT59), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n728_), .A2(new_n559_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n680_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n731_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n741_), .B2(new_n732_), .ZN(new_n742_));
  NOR4_X1   g541(.A1(new_n729_), .A2(KEYINPUT59), .A3(new_n731_), .A4(new_n733_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT119), .B(G113gat), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n411_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n737_), .B1(new_n744_), .B2(new_n746_), .ZN(G1340gat));
  INV_X1    g546(.A(G120gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n676_), .B2(KEYINPUT60), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n734_), .B(new_n749_), .C1(KEYINPUT60), .C2(new_n748_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n742_), .A2(new_n743_), .A3(new_n676_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT120), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT120), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n750_), .C1(new_n751_), .C2(new_n748_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1341gat));
  AOI21_X1  g555(.A(G127gat), .B1(new_n734_), .B2(new_n554_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n554_), .A2(G127gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n744_), .B2(new_n758_), .ZN(G1342gat));
  AOI21_X1  g558(.A(G134gat), .B1(new_n734_), .B2(new_n537_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n592_), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT121), .B(G134gat), .Z(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n744_), .B2(new_n763_), .ZN(G1343gat));
  INV_X1    g563(.A(new_n729_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n369_), .A2(new_n364_), .A3(new_n358_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n572_), .A3(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n411_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT122), .B(G141gat), .Z(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(new_n769_), .ZN(G1344gat));
  NOR2_X1   g569(.A1(new_n767_), .A2(new_n676_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(G148gat), .Z(G1345gat));
  OR3_X1    g571(.A1(new_n767_), .A2(KEYINPUT123), .A3(new_n559_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT123), .B1(new_n767_), .B2(new_n559_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(KEYINPUT61), .B(G155gat), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1346gat));
  INV_X1    g577(.A(G162gat), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n767_), .A2(new_n779_), .A3(new_n761_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n767_), .B2(new_n541_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT124), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n782_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(G1347gat));
  NOR2_X1   g584(.A1(new_n729_), .A2(new_n564_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n368_), .A2(new_n360_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n204_), .B1(new_n789_), .B2(new_n410_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT125), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(KEYINPUT62), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n786_), .A2(KEYINPUT126), .A3(new_n787_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT126), .B1(new_n786_), .B2(new_n787_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n243_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n410_), .A3(new_n796_), .ZN(new_n797_));
  XOR2_X1   g596(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n798_));
  OAI211_X1 g597(.A(new_n792_), .B(new_n797_), .C1(new_n790_), .C2(new_n798_), .ZN(G1348gat));
  OAI21_X1  g598(.A(G176gat), .B1(new_n788_), .B2(new_n676_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n795_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n507_), .A2(new_n205_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(G1349gat));
  AOI21_X1  g602(.A(G183gat), .B1(new_n789_), .B2(new_n554_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n559_), .A2(new_n209_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n795_), .B2(new_n805_), .ZN(G1350gat));
  OAI21_X1  g605(.A(G190gat), .B1(new_n801_), .B2(new_n761_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n795_), .A2(new_n537_), .A3(new_n210_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1351gat));
  NOR2_X1   g608(.A1(new_n242_), .A2(new_n322_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n765_), .A2(new_n360_), .A3(new_n369_), .A4(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n411_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n676_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g614(.A1(new_n811_), .A2(new_n559_), .ZN(new_n816_));
  OR2_X1    g615(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT127), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n816_), .A2(new_n817_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT127), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n816_), .A2(new_n822_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n820_), .A2(new_n821_), .A3(new_n823_), .ZN(G1354gat));
  NOR2_X1   g623(.A1(new_n811_), .A2(new_n541_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(G218gat), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n811_), .A2(new_n761_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(G218gat), .B2(new_n827_), .ZN(G1355gat));
endmodule


