//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_;
  NAND3_X1  g000(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT3), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT87), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT86), .B(KEYINPUT2), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  AND2_X1   g007(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n205_), .B(new_n207_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n202_), .B(new_n204_), .C1(new_n208_), .C2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(G155gat), .ZN(new_n215_));
  INV_X1    g014(.A(G162gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT29), .ZN(new_n219_));
  INV_X1    g018(.A(new_n203_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(KEYINPUT1), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT85), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT85), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n217_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n214_), .A2(KEYINPUT1), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n220_), .B(new_n207_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(new_n219_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  XNOR2_X1  g028(.A(G22gat), .B(G50gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G78gat), .B(G106gat), .Z(new_n233_));
  INV_X1    g032(.A(KEYINPUT93), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT89), .B(G204gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G197gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT21), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n240_), .A2(G204gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n235_), .B2(G197gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n238_), .B(new_n239_), .C1(new_n237_), .C2(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n240_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G197gat), .A2(G204gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(KEYINPUT21), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT90), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n246_), .A2(new_n250_), .A3(KEYINPUT21), .A4(new_n247_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G211gat), .B(G218gat), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n243_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n238_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n253_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n255_), .A2(KEYINPUT92), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT92), .B1(new_n255_), .B2(new_n257_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n219_), .B1(new_n218_), .B2(new_n226_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G228gat), .ZN(new_n262_));
  INV_X1    g061(.A(G233gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n234_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n255_), .A2(new_n257_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT92), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n260_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n255_), .A2(KEYINPUT92), .A3(new_n257_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT93), .A3(new_n264_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n233_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n233_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n275_), .ZN(new_n278_));
  AOI211_X1 g077(.A(new_n277_), .B(new_n278_), .C1(new_n266_), .C2(new_n273_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n232_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n274_), .A2(new_n233_), .A3(new_n275_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT95), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n272_), .A2(KEYINPUT93), .A3(new_n264_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT93), .B1(new_n272_), .B2(new_n264_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n275_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n277_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n274_), .A2(KEYINPUT95), .A3(new_n233_), .A4(new_n275_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n285_), .A2(new_n289_), .A3(new_n290_), .A4(new_n231_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n283_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(KEYINPUT94), .A3(new_n232_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n282_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n297_), .B(KEYINPUT82), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT82), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n298_), .A2(new_n299_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(new_n296_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT23), .ZN(new_n312_));
  OR3_X1    g111(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n304_), .A2(KEYINPUT83), .A3(new_n307_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G183gat), .ZN(new_n317_));
  INV_X1    g116(.A(G190gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G169gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n295_), .B1(new_n324_), .B2(new_n267_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(KEYINPUT96), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT96), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n312_), .A2(new_n327_), .A3(new_n319_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n322_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n302_), .A2(new_n296_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n314_), .A2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n325_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G64gat), .ZN(new_n343_));
  INV_X1    g142(.A(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n316_), .A2(new_n255_), .A3(new_n257_), .A4(new_n323_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n330_), .A2(new_n333_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n267_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(new_n349_), .A3(KEYINPUT20), .A4(new_n338_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n346_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n338_), .B1(new_n325_), .B2(new_n335_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n350_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n345_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT97), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n340_), .A2(new_n350_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(KEYINPUT97), .A3(new_n345_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n334_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n339_), .B1(new_n363_), .B2(new_n325_), .ZN(new_n364_));
  AND4_X1   g163(.A1(KEYINPUT20), .A2(new_n347_), .A3(new_n349_), .A4(new_n339_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n346_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT101), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n367_), .A2(new_n368_), .B1(new_n345_), .B2(new_n357_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n366_), .B2(KEYINPUT101), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n362_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(G127gat), .B(G134gat), .Z(new_n375_));
  INV_X1    g174(.A(G113gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G113gat), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n377_), .A2(G120gat), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(G120gat), .B1(new_n377_), .B2(new_n379_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n218_), .A2(new_n382_), .A3(new_n226_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n218_), .B2(new_n226_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n374_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n218_), .A2(new_n226_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n382_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT99), .B(KEYINPUT4), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n383_), .A2(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(KEYINPUT98), .A3(KEYINPUT4), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n218_), .A2(new_n382_), .A3(new_n226_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT98), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n390_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n385_), .B1(new_n397_), .B2(new_n374_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G85gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT0), .ZN(new_n401_));
  INV_X1    g200(.A(G57gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n405_), .B(new_n385_), .C1(new_n397_), .C2(new_n374_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n324_), .A2(KEYINPUT30), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n316_), .A2(new_n411_), .A3(new_n323_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT31), .B1(new_n413_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n413_), .A2(KEYINPUT31), .A3(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n382_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n420_), .A3(new_n387_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n410_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n423_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n408_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n294_), .A2(new_n373_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n404_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n390_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT98), .B1(new_n391_), .B2(KEYINPUT4), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n394_), .A2(new_n395_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n374_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT100), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT100), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n397_), .A2(new_n440_), .A3(new_n374_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n391_), .A2(new_n438_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n439_), .A2(new_n405_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n398_), .A2(KEYINPUT33), .A3(new_n403_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n433_), .A2(new_n443_), .A3(new_n359_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n357_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT32), .B(new_n345_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n407_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT94), .B1(new_n292_), .B2(new_n232_), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n281_), .B(new_n231_), .C1(new_n289_), .C2(new_n283_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n453_), .A3(new_n291_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n360_), .A2(new_n361_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n294_), .A2(new_n408_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n428_), .A2(new_n429_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n431_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G141gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT80), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G169gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(new_n240_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G29gat), .B(G36gat), .ZN(new_n464_));
  INV_X1    g263(.A(G43gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G50gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G8gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT76), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(G15gat), .A2(G22gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G15gat), .A2(G22gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G1gat), .A2(G8gat), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n472_), .A2(new_n473_), .B1(KEYINPUT14), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n471_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n468_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT79), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n468_), .B(KEYINPUT15), .ZN(new_n479_));
  INV_X1    g278(.A(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n468_), .A2(new_n476_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n482_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n463_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n463_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n478_), .A2(new_n485_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n483_), .B(new_n488_), .C1(new_n489_), .C2(new_n482_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(KEYINPUT81), .B(new_n463_), .C1(new_n484_), .C2(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G148gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G176gat), .B(G204gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT73), .B(G120gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G57gat), .B(G64gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n503_), .A2(KEYINPUT11), .ZN(new_n504_));
  XOR2_X1   g303(.A(G71gat), .B(G78gat), .Z(new_n505_));
  OR2_X1    g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n503_), .A2(KEYINPUT11), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n505_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n509_), .A2(KEYINPUT12), .ZN(new_n510_));
  INV_X1    g309(.A(G85gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT65), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT65), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G85gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n514_), .A3(G92gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT66), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n519_));
  AND3_X1   g318(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT67), .B1(new_n511_), .B2(new_n344_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n522_), .B1(new_n523_), .B2(new_n520_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n518_), .A2(new_n519_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(G99gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT10), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT10), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G99gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT64), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n526_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT6), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(new_n538_), .A3(KEYINPUT68), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT68), .B1(new_n536_), .B2(new_n538_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT69), .B1(new_n525_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n528_), .A2(new_n530_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT64), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n546_));
  AOI21_X1  g345(.A(G106gat), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n537_), .B1(G99gat), .B2(G106gat), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n535_), .A2(KEYINPUT6), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n536_), .A2(new_n538_), .A3(KEYINPUT68), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n515_), .A2(new_n517_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT66), .ZN(new_n556_));
  NAND3_X1  g355(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n557_));
  MUX2_X1   g356(.A(KEYINPUT67), .B(new_n523_), .S(new_n557_), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n554_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n543_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n564_));
  OR3_X1    g363(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n551_), .A2(new_n552_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G85gat), .B(G92gat), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT8), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n549_), .A2(new_n550_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n564_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n567_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n566_), .A2(new_n569_), .B1(new_n572_), .B2(KEYINPUT8), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT71), .B1(new_n563_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n576_), .B(new_n573_), .C1(new_n543_), .C2(new_n562_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n510_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n509_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n525_), .A2(new_n542_), .A3(KEYINPUT69), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n561_), .B1(new_n554_), .B2(new_n560_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n574_), .B(new_n579_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT12), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n574_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n509_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n578_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n582_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(G230gat), .A3(G233gat), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n502_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n502_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n501_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n591_), .A2(new_n592_), .A3(new_n501_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n598_));
  OAI22_X1  g397(.A1(new_n594_), .A2(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n595_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n459_), .A2(new_n494_), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n563_), .A2(new_n468_), .A3(new_n574_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT75), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n479_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n606_), .B(new_n607_), .C1(KEYINPUT35), .C2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(G134gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n216_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n606_), .A2(KEYINPUT35), .A3(new_n609_), .A4(new_n607_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n612_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n612_), .A2(new_n618_), .B1(new_n616_), .B2(new_n615_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n612_), .A2(new_n618_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n615_), .A2(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n612_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT37), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n509_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n476_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT17), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT17), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n632_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n638_), .B2(new_n632_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT78), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n623_), .A2(new_n629_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n604_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n644_), .A2(G1gat), .A3(new_n408_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT103), .B1(new_n459_), .B2(new_n628_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n603_), .A2(new_n494_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649_));
  INV_X1    g448(.A(new_n458_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n649_), .B(new_n621_), .C1(new_n651_), .C2(new_n431_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n647_), .A2(new_n648_), .A3(new_n642_), .A4(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n408_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n646_), .A2(new_n654_), .A3(new_n655_), .ZN(G1324gat));
  OAI21_X1  g455(.A(G8gat), .B1(new_n653_), .B2(new_n455_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n659_), .B(G8gat), .C1(new_n653_), .C2(new_n455_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n455_), .A2(G8gat), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n644_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT104), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(new_n667_), .A3(new_n664_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT40), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT104), .B(new_n663_), .C1(new_n658_), .C2(new_n660_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n669_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n653_), .B2(new_n458_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT41), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n644_), .A2(G15gat), .A3(new_n458_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(new_n294_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n644_), .A2(G22gat), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n653_), .B2(new_n679_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT105), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT105), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(KEYINPUT42), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT42), .B1(new_n682_), .B2(new_n683_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(G29gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n623_), .A2(new_n629_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n459_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n691_), .B(new_n688_), .C1(new_n651_), .C2(new_n431_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n642_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n648_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n648_), .A4(new_n694_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n687_), .B1(new_n699_), .B2(new_n407_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n621_), .A2(new_n642_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n604_), .A2(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(G29gat), .A3(new_n408_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1328gat));
  NOR3_X1   g503(.A1(new_n702_), .A2(G36gat), .A3(new_n455_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT45), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n373_), .A3(new_n698_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n707_), .B2(G36gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI221_X1 g511(.A(new_n706_), .B1(KEYINPUT107), .B2(KEYINPUT46), .C1(new_n708_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  AOI21_X1  g513(.A(new_n465_), .B1(new_n699_), .B2(new_n650_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n702_), .A2(G43gat), .A3(new_n458_), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n697_), .A2(new_n294_), .A3(new_n698_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n697_), .A2(KEYINPUT108), .A3(new_n294_), .A4(new_n698_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(G50gat), .A3(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n604_), .A2(new_n467_), .A3(new_n294_), .A4(new_n701_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT109), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n725_), .A2(new_n729_), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1331gat));
  INV_X1    g530(.A(new_n494_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n602_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n647_), .A2(new_n642_), .A3(new_n652_), .A4(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n408_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n733_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n459_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n643_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n407_), .A2(new_n402_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT110), .Z(G1332gat));
  OAI21_X1  g540(.A(G64gat), .B1(new_n734_), .B2(new_n455_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n455_), .A2(G64gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n738_), .B2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n734_), .B2(new_n458_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n458_), .A2(G71gat), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT111), .Z(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n738_), .B2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n734_), .B2(new_n679_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT50), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n679_), .A2(G78gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n738_), .B2(new_n753_), .ZN(G1335gat));
  AOI21_X1  g553(.A(new_n736_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n694_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n756_), .A2(new_n407_), .A3(new_n512_), .A4(new_n514_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n737_), .A2(new_n701_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n511_), .B1(new_n758_), .B2(new_n408_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT112), .Z(G1336gat));
  NOR3_X1   g560(.A1(new_n758_), .A2(G92gat), .A3(new_n455_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n756_), .A2(new_n373_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G92gat), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT113), .ZN(G1337gat));
  AOI211_X1 g564(.A(new_n458_), .B(new_n758_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n756_), .A2(new_n650_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G99gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g568(.A1(new_n693_), .A2(new_n694_), .A3(new_n294_), .A4(new_n733_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n755_), .A2(KEYINPUT114), .A3(new_n694_), .A4(new_n294_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(G106gat), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT52), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n772_), .A2(new_n776_), .A3(G106gat), .A4(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n737_), .A2(new_n526_), .A3(new_n294_), .A4(new_n701_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n782_), .A3(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  INV_X1    g583(.A(new_n482_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n478_), .A2(new_n481_), .A3(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n463_), .B(new_n786_), .C1(new_n489_), .C2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n490_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n600_), .B2(new_n593_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n587_), .B1(new_n578_), .B2(new_n586_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n588_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n578_), .A2(new_n586_), .A3(KEYINPUT55), .A4(new_n587_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n790_), .B1(new_n795_), .B2(new_n501_), .ZN(new_n796_));
  AOI211_X1 g595(.A(KEYINPUT56), .B(new_n500_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n595_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n789_), .B1(new_n798_), .B2(new_n732_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT115), .B1(new_n799_), .B2(new_n628_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(new_n796_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n795_), .A2(new_n790_), .A3(new_n501_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(new_n732_), .A3(new_n600_), .A4(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n789_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n621_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(new_n801_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(KEYINPUT57), .A3(new_n621_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n788_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n802_), .A2(new_n600_), .A3(new_n811_), .A4(new_n803_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT116), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT58), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT116), .A3(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n688_), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n809_), .A2(new_n810_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n694_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n643_), .A2(new_n602_), .A3(new_n820_), .A4(new_n494_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n623_), .A2(new_n629_), .A3(new_n494_), .A4(new_n642_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n822_), .B2(new_n603_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n824_), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n294_), .A2(new_n373_), .A3(new_n458_), .A4(new_n408_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n732_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n824_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n809_), .A2(new_n817_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n809_), .A2(KEYINPUT117), .A3(new_n817_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n810_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n830_), .B1(new_n835_), .B2(new_n694_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n826_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n837_), .A2(new_n840_), .B1(KEYINPUT59), .B2(new_n827_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n494_), .A2(new_n376_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n829_), .B1(new_n841_), .B2(new_n842_), .ZN(G1340gat));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n602_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n828_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n603_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n848_), .B2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g648(.A(G127gat), .B1(new_n828_), .B2(new_n642_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n642_), .A2(G127gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n841_), .B2(new_n851_), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(new_n828_), .B2(new_n628_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n688_), .A2(G134gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n841_), .B2(new_n854_), .ZN(G1343gat));
  AOI21_X1  g654(.A(new_n830_), .B1(new_n818_), .B2(new_n694_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n679_), .A2(new_n373_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n407_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n856_), .A2(new_n650_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n732_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n603_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g662(.A(new_n858_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n825_), .A2(new_n642_), .A3(new_n458_), .A4(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT118), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n856_), .A2(new_n650_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n868_), .A2(new_n869_), .A3(new_n642_), .A4(new_n864_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n866_), .A2(new_n867_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n866_), .B2(new_n870_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n215_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n865_), .A2(KEYINPUT118), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n869_), .B1(new_n859_), .B2(new_n642_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT61), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n866_), .A2(new_n867_), .A3(new_n870_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G155gat), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n873_), .A2(new_n878_), .ZN(G1346gat));
  AOI21_X1  g678(.A(G162gat), .B1(new_n859_), .B2(new_n628_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n689_), .A2(new_n216_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n859_), .B2(new_n881_), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n430_), .A2(new_n455_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT119), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n679_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n836_), .A2(new_n494_), .A3(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n298_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT120), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n888_), .A2(KEYINPUT120), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n298_), .A2(KEYINPUT22), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n298_), .A2(KEYINPUT22), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n886_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT120), .B(new_n888_), .C1(new_n886_), .C2(new_n298_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n894_), .A3(new_n895_), .ZN(G1348gat));
  NOR2_X1   g695(.A1(new_n836_), .A2(new_n885_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G176gat), .B1(new_n897_), .B2(new_n603_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n856_), .A2(new_n294_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n899_), .A2(G176gat), .A3(new_n884_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n603_), .B2(new_n900_), .ZN(G1349gat));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n642_), .A3(new_n884_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n903_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n317_), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n305_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n897_), .A2(new_n642_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT121), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n897_), .A2(new_n910_), .A3(new_n642_), .A4(new_n907_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n906_), .A2(new_n909_), .A3(new_n911_), .ZN(G1350gat));
  NAND2_X1  g711(.A1(new_n628_), .A2(new_n306_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT123), .Z(new_n914_));
  NAND2_X1  g713(.A1(new_n897_), .A2(new_n914_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n836_), .A2(new_n689_), .A3(new_n885_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n318_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n294_), .A2(new_n408_), .A3(new_n458_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n455_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n825_), .A2(new_n732_), .A3(new_n920_), .A4(new_n921_), .ZN(new_n922_));
  OR3_X1    g721(.A1(new_n922_), .A2(KEYINPUT126), .A3(new_n240_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT126), .B1(new_n922_), .B2(new_n240_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT125), .B1(new_n922_), .B2(new_n240_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n825_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n602_), .ZN(new_n929_));
  MUX2_X1   g728(.A(G204gat), .B(new_n235_), .S(new_n929_), .Z(G1353gat));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n694_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AND2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  NOR2_X1   g734(.A1(new_n928_), .A2(new_n621_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n688_), .A2(G218gat), .ZN(new_n937_));
  OAI22_X1  g736(.A1(new_n936_), .A2(G218gat), .B1(new_n928_), .B2(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


