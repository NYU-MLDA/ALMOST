//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT7), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n202_), .A2(new_n212_), .A3(new_n203_), .A4(new_n204_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n206_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n221_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n214_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n214_), .B2(new_n220_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n204_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT10), .B(G99gat), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n233_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n227_), .B(new_n229_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G78gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(G57gat), .B(G64gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(KEYINPUT11), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n237_), .B2(KEYINPUT11), .ZN(new_n240_));
  INV_X1    g039(.A(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G57gat), .ZN(new_n242_));
  INV_X1    g041(.A(G57gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G64gat), .ZN(new_n244_));
  AND4_X1   g043(.A1(new_n239_), .A2(new_n242_), .A3(new_n244_), .A4(KEYINPUT11), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n238_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n244_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n237_), .A2(new_n239_), .A3(KEYINPUT11), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n248_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .A4(new_n236_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n246_), .A2(new_n252_), .A3(KEYINPUT68), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT68), .B1(new_n246_), .B2(new_n252_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n226_), .B(new_n235_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n246_), .A2(new_n252_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n214_), .A2(new_n220_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n223_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n214_), .A2(new_n223_), .A3(new_n220_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n235_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n246_), .A2(new_n252_), .A3(KEYINPUT68), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G230gat), .A2(G233gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n255_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n255_), .B2(new_n267_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n224_), .A2(new_n225_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT69), .B1(new_n261_), .B2(new_n262_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n235_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n256_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT12), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(KEYINPUT70), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282_));
  INV_X1    g081(.A(new_n235_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n274_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n261_), .A2(KEYINPUT69), .A3(new_n262_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n286_), .B2(new_n279_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT12), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n265_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n269_), .B1(new_n273_), .B2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G120gat), .B(G148gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(G176gat), .B(G204gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n269_), .B(new_n296_), .C1(new_n273_), .C2(new_n290_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G29gat), .B(G36gat), .Z(new_n305_));
  XOR2_X1   g104(.A(G43gat), .B(G50gat), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G29gat), .B(G36gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G43gat), .B(G50gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT15), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  INV_X1    g112(.A(G1gat), .ZN(new_n314_));
  INV_X1    g113(.A(G8gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT14), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G1gat), .B(G8gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n311_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G229gat), .A2(G233gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT76), .Z(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n319_), .B(new_n321_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(G229gat), .A3(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G113gat), .B(G141gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G169gat), .B(G197gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT77), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n325_), .A2(new_n327_), .A3(new_n333_), .A4(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n325_), .A2(new_n327_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n304_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT90), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  OR2_X1    g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  OR3_X1    g143(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT84), .ZN(new_n347_));
  INV_X1    g146(.A(G141gat), .ZN(new_n348_));
  INV_X1    g147(.A(G148gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n345_), .B(new_n346_), .C1(new_n350_), .C2(KEYINPUT2), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(KEYINPUT2), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n343_), .B(new_n344_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n343_), .A2(KEYINPUT1), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G155gat), .A3(G162gat), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n354_), .A2(new_n356_), .A3(new_n344_), .A4(KEYINPUT83), .ZN(new_n357_));
  XOR2_X1   g156(.A(G141gat), .B(G148gat), .Z(new_n358_));
  OAI211_X1 g157(.A(new_n357_), .B(new_n358_), .C1(KEYINPUT83), .C2(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT85), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT21), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT86), .B(G204gat), .ZN(new_n364_));
  INV_X1    g163(.A(G197gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n367_));
  INV_X1    g166(.A(G204gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(G197gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n364_), .A2(new_n367_), .A3(new_n365_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n363_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G211gat), .B(G218gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n364_), .A2(G197gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n363_), .B1(G197gat), .B2(G204gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n370_), .A2(new_n371_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n373_), .A2(new_n363_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n360_), .A2(new_n383_), .A3(KEYINPUT29), .ZN(new_n384_));
  INV_X1    g183(.A(G228gat), .ZN(new_n385_));
  INV_X1    g184(.A(G233gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n362_), .A2(new_n382_), .A3(new_n384_), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n372_), .A2(new_n377_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(new_n387_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n393_), .A2(KEYINPUT88), .A3(new_n384_), .A4(new_n362_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n388_), .B1(new_n382_), .B2(new_n361_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n341_), .B(new_n342_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n342_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT90), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n342_), .B(KEYINPUT89), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT28), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G22gat), .B(G50gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n397_), .A2(new_n400_), .A3(new_n402_), .A4(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n402_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n398_), .A2(new_n401_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n360_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G127gat), .B(G134gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G113gat), .B(G120gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT82), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n414_), .A2(new_n415_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n360_), .B1(new_n418_), .B2(new_n416_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT4), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n360_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n421_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n423_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n429_), .A2(new_n437_), .A3(new_n432_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n443_));
  NOR2_X1   g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G169gat), .ZN(new_n447_));
  INV_X1    g246(.A(G176gat), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n446_), .B(KEYINPUT24), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT25), .B(G183gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT78), .ZN(new_n454_));
  INV_X1    g253(.A(G190gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT26), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n455_), .A2(KEYINPUT26), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n453_), .B(new_n456_), .C1(new_n457_), .C2(new_n454_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n444_), .B(KEYINPUT79), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT24), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n449_), .A2(new_n452_), .A3(new_n458_), .A4(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G183gat), .A2(G190gat), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n450_), .A2(new_n451_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n466_));
  OR3_X1    g265(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT80), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n471_), .A3(new_n468_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n392_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT26), .B(G190gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n453_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n444_), .A2(new_n460_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n476_), .A2(new_n452_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n449_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT22), .B(G169gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT92), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(G176gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n447_), .A2(new_n448_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n464_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n479_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n474_), .B1(new_n382_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n473_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G226gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n392_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n491_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT20), .B(new_n494_), .C1(new_n382_), .C2(new_n486_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT93), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n472_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n471_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n382_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n486_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n474_), .B1(new_n500_), .B2(new_n392_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT93), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(new_n501_), .A3(new_n502_), .A4(new_n494_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n492_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT18), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G64gat), .B(G92gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n492_), .A2(new_n496_), .A3(new_n503_), .A4(new_n508_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n443_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n488_), .A2(new_n491_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n501_), .A2(KEYINPUT94), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT20), .B1(new_n382_), .B2(new_n486_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n518_), .A3(new_n499_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n491_), .B2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(KEYINPUT27), .B(new_n511_), .C1(new_n520_), .C2(new_n508_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n412_), .A2(new_n442_), .A3(new_n513_), .A4(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n508_), .A2(KEYINPUT32), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n492_), .A2(new_n496_), .A3(new_n503_), .A4(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n441_), .B(new_n524_), .C1(new_n520_), .C2(new_n523_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n437_), .B1(new_n431_), .B2(new_n423_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n424_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT33), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n439_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n433_), .A2(KEYINPUT33), .A3(new_n438_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n529_), .A2(new_n510_), .A3(new_n511_), .A4(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n411_), .A3(new_n407_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n522_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n419_), .B(KEYINPUT31), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G99gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G15gat), .B(G43gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT81), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT30), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n470_), .A2(new_n472_), .A3(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(G71gat), .Z(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n546_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n537_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n547_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n536_), .A3(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n534_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n521_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT96), .B1(new_n556_), .B2(new_n512_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n513_), .A2(new_n558_), .A3(new_n521_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n412_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n442_), .A3(new_n561_), .A4(new_n553_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n340_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n566_));
  INV_X1    g365(.A(new_n312_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n286_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n263_), .A2(new_n321_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n566_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(new_n569_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n566_), .A2(new_n573_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n570_), .A2(new_n571_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n570_), .A2(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G134gat), .B(G162gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(new_n581_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n575_), .A2(new_n576_), .A3(new_n581_), .A4(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(KEYINPUT37), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n258_), .A2(new_n264_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT75), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n319_), .B(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n596_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n600_), .A2(new_n278_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n603_), .A2(new_n595_), .A3(new_n594_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n278_), .B2(new_n600_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n590_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n563_), .A2(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT97), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT97), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n609_), .A2(new_n314_), .A3(new_n441_), .A4(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n612_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n586_), .B(KEYINPUT98), .Z(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n606_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n563_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n442_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(new_n614_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n613_), .A2(KEYINPUT99), .A3(new_n614_), .A4(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1324gat));
  NOR3_X1   g422(.A1(new_n556_), .A2(KEYINPUT96), .A3(new_n512_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n558_), .B1(new_n513_), .B2(new_n521_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n563_), .A2(new_n626_), .A3(new_n616_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G8gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT39), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n609_), .A2(new_n315_), .A3(new_n626_), .A4(new_n610_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n617_), .B2(new_n554_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n554_), .A2(G15gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n608_), .B2(new_n637_), .ZN(G1326gat));
  XOR2_X1   g437(.A(new_n412_), .B(KEYINPUT102), .Z(new_n639_));
  OR3_X1    g438(.A1(new_n608_), .A2(G22gat), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G22gat), .B1(new_n617_), .B2(new_n639_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT42), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(KEYINPUT42), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT103), .Z(G1327gat));
  INV_X1    g444(.A(G29gat), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  INV_X1    g446(.A(new_n590_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n649_), .B2(KEYINPUT105), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n407_), .A2(new_n553_), .A3(new_n411_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n441_), .B(new_n651_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n553_), .B1(new_n522_), .B2(new_n533_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n590_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(KEYINPUT43), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n606_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n340_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT104), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT104), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT44), .B1(new_n657_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n665_), .B(new_n662_), .C1(new_n650_), .C2(new_n656_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n646_), .B1(new_n667_), .B2(new_n441_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n586_), .A2(new_n658_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n563_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n441_), .A2(new_n646_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT106), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT107), .B1(new_n668_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n664_), .A2(new_n666_), .A3(new_n442_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n677_), .B(new_n674_), .C1(new_n678_), .C2(new_n646_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  INV_X1    g480(.A(G36gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n667_), .B2(new_n626_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n626_), .A2(KEYINPUT108), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n626_), .A2(KEYINPUT108), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n682_), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n687_), .A2(KEYINPUT45), .A3(new_n670_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT45), .B1(new_n687_), .B2(new_n670_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n681_), .B1(new_n683_), .B2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n664_), .A2(new_n666_), .A3(new_n560_), .ZN(new_n693_));
  OAI211_X1 g492(.A(KEYINPUT46), .B(new_n690_), .C1(new_n693_), .C2(new_n682_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(G43gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n554_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n667_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n670_), .B2(new_n554_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n702_), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1330gat));
  INV_X1    g503(.A(new_n639_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G50gat), .B1(new_n671_), .B2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n412_), .A2(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n667_), .B2(new_n707_), .ZN(G1331gat));
  NAND2_X1  g507(.A1(new_n555_), .A2(new_n562_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n304_), .A2(new_n339_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n616_), .A3(new_n710_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(KEYINPUT111), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(KEYINPUT111), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n714_), .A2(new_n243_), .A3(new_n442_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n709_), .A2(new_n710_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n607_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n442_), .B1(new_n717_), .B2(KEYINPUT109), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(KEYINPUT109), .B2(new_n717_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n243_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(KEYINPUT110), .A3(new_n243_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n715_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(new_n717_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n241_), .A3(new_n686_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n712_), .A2(new_n686_), .A3(new_n713_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(G64gat), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G64gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT113), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n726_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1333gat));
  OR3_X1    g534(.A1(new_n717_), .A2(G71gat), .A3(new_n554_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n714_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n553_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT49), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G71gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G71gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(G1334gat));
  INV_X1    g541(.A(G78gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n725_), .A2(new_n743_), .A3(new_n705_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n737_), .B2(new_n705_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n710_), .A2(new_n606_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n650_), .B2(new_n656_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n442_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n716_), .A2(new_n669_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n215_), .A3(new_n441_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(G1336gat));
  INV_X1    g556(.A(new_n686_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G92gat), .B1(new_n752_), .B2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n216_), .A3(new_n626_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1337gat));
  NOR3_X1   g560(.A1(new_n754_), .A2(new_n233_), .A3(new_n554_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n751_), .A2(new_n553_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G99gat), .ZN(new_n764_));
  NAND2_X1  g563(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(G1338gat));
  AOI21_X1  g565(.A(new_n204_), .B1(KEYINPUT116), .B2(KEYINPUT52), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n751_), .B2(new_n412_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n755_), .A2(new_n204_), .A3(new_n412_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT53), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n769_), .A2(new_n771_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(G1339gat));
  INV_X1    g579(.A(new_n339_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n304_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n339_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n607_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n607_), .B2(new_n783_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n339_), .A2(new_n299_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT117), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n339_), .A2(new_n790_), .A3(new_n299_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n273_), .B2(new_n290_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n281_), .A2(new_n287_), .A3(new_n255_), .A4(new_n289_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n268_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n263_), .B1(new_n258_), .B2(new_n264_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT71), .B1(new_n798_), .B2(new_n268_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n255_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n284_), .A2(new_n285_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n279_), .B1(new_n802_), .B2(new_n235_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n803_), .A2(KEYINPUT70), .B1(new_n288_), .B2(new_n265_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n801_), .A2(new_n804_), .A3(KEYINPUT55), .A4(new_n287_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n794_), .A2(new_n797_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n796_), .B1(new_n795_), .B2(new_n268_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n297_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT56), .B(new_n297_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n792_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n330_), .B1(new_n326_), .B2(new_n324_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n320_), .A2(new_n322_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n324_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n335_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n300_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n586_), .B1(new_n812_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT57), .B(new_n586_), .C1(new_n812_), .C2(new_n818_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n816_), .A2(new_n299_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n823_), .B(new_n590_), .C1(new_n825_), .C2(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n824_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n811_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n795_), .A2(new_n268_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT118), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(new_n797_), .A3(new_n794_), .A4(new_n805_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n297_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n829_), .B1(new_n830_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n823_), .B1(new_n837_), .B2(new_n590_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n821_), .B(new_n822_), .C1(new_n828_), .C2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n787_), .B1(new_n839_), .B2(new_n606_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n442_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n626_), .A2(new_n651_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(KEYINPUT59), .A3(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n821_), .A2(new_n822_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n590_), .B1(new_n825_), .B2(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT119), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n658_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n441_), .B(new_n842_), .C1(new_n848_), .C2(new_n787_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n781_), .B1(new_n843_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G113gat), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n339_), .A2(new_n853_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n852_), .A2(new_n853_), .B1(new_n849_), .B2(new_n854_), .ZN(G1340gat));
  AOI21_X1  g654(.A(new_n304_), .B1(new_n843_), .B2(new_n851_), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n304_), .B2(KEYINPUT60), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(KEYINPUT60), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(KEYINPUT120), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(KEYINPUT120), .B2(new_n858_), .ZN(new_n861_));
  OAI22_X1  g660(.A1(new_n856_), .A2(new_n857_), .B1(new_n849_), .B2(new_n861_), .ZN(G1341gat));
  AOI21_X1  g661(.A(new_n606_), .B1(new_n843_), .B2(new_n851_), .ZN(new_n863_));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n658_), .A2(new_n864_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n863_), .A2(new_n864_), .B1(new_n849_), .B2(new_n865_), .ZN(G1342gat));
  NAND3_X1  g665(.A1(new_n841_), .A2(new_n842_), .A3(new_n615_), .ZN(new_n867_));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT121), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n590_), .A2(G134gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n843_), .B2(new_n851_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n615_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT121), .B(new_n868_), .C1(new_n849_), .C2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n869_), .A2(new_n871_), .A3(new_n874_), .ZN(G1343gat));
  NOR3_X1   g674(.A1(new_n686_), .A2(new_n561_), .A3(new_n553_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n841_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n781_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n348_), .ZN(G1344gat));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n304_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n349_), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n841_), .A2(new_n658_), .A3(new_n876_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n877_), .B2(new_n648_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n872_), .A2(G162gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n877_), .B2(new_n886_), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n554_), .A2(new_n441_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n686_), .A2(new_n639_), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n840_), .B2(new_n890_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n686_), .A2(new_n639_), .A3(new_n889_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT122), .B(new_n892_), .C1(new_n848_), .C2(new_n787_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n481_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n339_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n840_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(new_n339_), .A3(new_n892_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n896_), .B1(new_n900_), .B2(new_n901_), .ZN(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n894_), .B2(new_n782_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n897_), .A2(new_n561_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n686_), .A2(new_n889_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(G176gat), .A3(new_n782_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT123), .B1(new_n903_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n304_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n910_));
  OAI221_X1 g709(.A(new_n909_), .B1(new_n904_), .B2(new_n906_), .C1(new_n910_), .C2(G176gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n911_), .ZN(G1349gat));
  NOR2_X1   g711(.A1(new_n606_), .A2(new_n453_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n897_), .A2(new_n561_), .A3(new_n658_), .A4(new_n905_), .ZN(new_n914_));
  INV_X1    g713(.A(G183gat), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n894_), .A2(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n894_), .A2(new_n475_), .A3(new_n615_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n648_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n455_), .ZN(G1351gat));
  NOR4_X1   g718(.A1(new_n758_), .A2(new_n441_), .A3(new_n561_), .A4(new_n553_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n897_), .A2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n339_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT124), .B(G197gat), .Z(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1352gat));
  NAND3_X1  g723(.A1(new_n897_), .A2(new_n920_), .A3(new_n782_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n368_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n897_), .A2(new_n920_), .A3(new_n782_), .A4(new_n364_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1353gat));
  NAND3_X1  g730(.A1(new_n897_), .A2(new_n920_), .A3(new_n658_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT63), .B(G211gat), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n897_), .A2(new_n920_), .A3(new_n658_), .A4(new_n935_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n933_), .A2(new_n934_), .A3(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n933_), .B2(new_n936_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1354gat));
  AOI21_X1  g738(.A(G218gat), .B1(new_n921_), .B2(new_n615_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n590_), .A2(G218gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n921_), .B2(new_n942_), .ZN(G1355gat));
endmodule


