//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G71gat), .B(G78gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT11), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n207_));
  INV_X1    g006(.A(new_n205_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n212_), .B(new_n213_), .C1(new_n215_), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n218_), .A2(KEYINPUT8), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT8), .B1(new_n218_), .B2(new_n224_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n215_), .A2(new_n217_), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT10), .B(G99gat), .Z(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n222_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n232_), .A2(new_n233_), .B1(KEYINPUT9), .B2(new_n220_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n234_), .B(new_n235_), .C1(KEYINPUT9), .C2(new_n223_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT9), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT9), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n221_), .A2(new_n222_), .B1(new_n238_), .B2(G92gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n231_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n211_), .B1(new_n227_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n203_), .B1(new_n242_), .B2(KEYINPUT12), .ZN(new_n243_));
  INV_X1    g042(.A(new_n226_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n218_), .A2(KEYINPUT8), .A3(new_n224_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n211_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT12), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT68), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(KEYINPUT12), .A3(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT67), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n242_), .A2(new_n254_), .A3(KEYINPUT12), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n241_), .A2(new_n244_), .A3(new_n245_), .A4(new_n211_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT69), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n251_), .A2(new_n256_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT70), .ZN(new_n267_));
  INV_X1    g066(.A(new_n260_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n257_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(new_n242_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n251_), .A2(new_n256_), .A3(new_n265_), .A4(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G120gat), .B(G148gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n267_), .A2(new_n270_), .A3(new_n272_), .A4(new_n278_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(KEYINPUT72), .A3(new_n279_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT13), .B1(new_n283_), .B2(new_n284_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n202_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n284_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT13), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT73), .A3(new_n285_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT74), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT107), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT99), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G197gat), .A2(G204gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G197gat), .A2(G204gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(KEYINPUT21), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  AND2_X1   g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(new_n299_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n302_), .A2(new_n305_), .A3(KEYINPUT95), .A4(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT95), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n307_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT25), .B(G183gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT26), .B(G190gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(G169gat), .B2(G176gat), .ZN(new_n315_));
  INV_X1    g114(.A(G169gat), .ZN(new_n316_));
  INV_X1    g115(.A(G176gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n312_), .A2(new_n313_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n316_), .A2(new_n317_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT22), .B(G169gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(new_n317_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n323_), .B(new_n324_), .C1(G183gat), .C2(G190gat), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n319_), .A2(new_n326_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n298_), .B1(new_n311_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n319_), .A2(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n336_), .B(new_n309_), .C1(new_n302_), .C2(new_n306_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(KEYINPUT99), .A4(new_n307_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n297_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G169gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n316_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(new_n317_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT86), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n344_), .B(new_n330_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n315_), .A2(new_n318_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G183gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n322_), .A2(KEYINPUT26), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT26), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G190gat), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .A4(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT83), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n346_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n357_), .A2(KEYINPUT84), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n326_), .B1(new_n357_), .B2(KEYINPUT84), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n345_), .B(new_n311_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n339_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT19), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n345_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n311_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n311_), .A2(new_n331_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT20), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT18), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND3_X1  g175(.A1(new_n364_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT105), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(KEYINPUT105), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT27), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n339_), .A2(new_n360_), .A3(new_n368_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n370_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n368_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n376_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(new_n379_), .A3(new_n385_), .ZN(new_n386_));
  AOI211_X1 g185(.A(new_n363_), .B(new_n370_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n368_), .B1(new_n339_), .B2(new_n360_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n384_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n377_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT106), .B1(new_n390_), .B2(new_n380_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT106), .ZN(new_n392_));
  AOI211_X1 g191(.A(new_n392_), .B(KEYINPUT27), .C1(new_n389_), .C2(new_n377_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n386_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT90), .B1(new_n395_), .B2(KEYINPUT1), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(G155gat), .A4(G162gat), .ZN(new_n399_));
  OR2_X1    g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(KEYINPUT1), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n396_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(KEYINPUT2), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(G141gat), .A3(G148gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n403_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n403_), .A2(new_n413_), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT91), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(new_n414_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n400_), .A2(new_n395_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n417_), .A2(KEYINPUT92), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT92), .B1(new_n417_), .B2(new_n418_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n407_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G127gat), .B(G134gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(G113gat), .B(G120gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n426_), .B(new_n407_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(KEYINPUT4), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(new_n431_), .A3(new_n424_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  NAND3_X1  g236(.A1(new_n425_), .A2(new_n429_), .A3(new_n427_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n433_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT104), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT104), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n439_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n407_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n417_), .A2(new_n418_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n417_), .A2(KEYINPUT92), .A3(new_n418_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n446_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT29), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n366_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(G228gat), .B(G233gat), .C1(new_n311_), .C2(KEYINPUT96), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n311_), .B1(new_n421_), .B2(KEYINPUT29), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT97), .Z(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n456_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G22gat), .B(G50gat), .Z(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n467_));
  OR3_X1    g266(.A1(new_n421_), .A2(KEYINPUT29), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n421_), .B2(KEYINPUT29), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n466_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT94), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n474_));
  INV_X1    g273(.A(new_n472_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(new_n470_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n465_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n475_), .A2(new_n470_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n461_), .A2(KEYINPUT98), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n459_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n459_), .A2(new_n479_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n442_), .B(new_n445_), .C1(new_n477_), .C2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n394_), .A2(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n389_), .A2(new_n377_), .A3(KEYINPUT100), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT100), .B1(new_n389_), .B2(new_n377_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n439_), .A2(KEYINPUT33), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n433_), .A2(new_n489_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT101), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n449_), .A2(new_n450_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n426_), .B1(new_n493_), .B2(new_n407_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n427_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n492_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n425_), .A2(KEYINPUT101), .A3(new_n427_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n430_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n437_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT102), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(KEYINPUT102), .A3(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n428_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n491_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT103), .B1(new_n487_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT100), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n387_), .A2(new_n388_), .A3(new_n384_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n376_), .B1(new_n364_), .B2(new_n372_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n389_), .A2(new_n377_), .A3(KEYINPUT100), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT103), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n498_), .A2(new_n499_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT102), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n502_), .A3(new_n501_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n511_), .A2(new_n512_), .A3(new_n516_), .A4(new_n491_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n387_), .A2(new_n388_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n376_), .A2(KEYINPUT32), .ZN(new_n519_));
  MUX2_X1   g318(.A(new_n383_), .B(new_n518_), .S(new_n519_), .Z(new_n520_));
  NOR2_X1   g319(.A1(new_n440_), .A2(new_n441_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n505_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n477_), .A2(new_n482_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n484_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G15gat), .B(G43gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G71gat), .B(G99gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n365_), .B(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(KEYINPUT87), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT30), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n530_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT89), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n535_), .A2(new_n536_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n424_), .B(KEYINPUT31), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n538_), .A2(new_n542_), .A3(new_n543_), .A4(new_n540_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n296_), .B1(new_n526_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n442_), .A2(new_n445_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT108), .ZN(new_n551_));
  INV_X1    g350(.A(new_n394_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n525_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n525_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n554_), .A2(new_n394_), .A3(KEYINPUT108), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n547_), .B(new_n550_), .C1(new_n553_), .C2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n545_), .A2(new_n546_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n516_), .B(new_n491_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n522_), .B1(new_n558_), .B2(KEYINPUT103), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n554_), .B1(new_n559_), .B2(new_n517_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT107), .B(new_n557_), .C1(new_n560_), .C2(new_n484_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n548_), .A2(new_n556_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563_));
  INV_X1    g362(.A(G1gat), .ZN(new_n564_));
  INV_X1    g363(.A(G8gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G1gat), .B(G8gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G29gat), .B(G36gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G43gat), .B(G50gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n569_), .B(new_n572_), .Z(new_n573_));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n572_), .B(KEYINPUT15), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n569_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n569_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n575_), .B1(new_n578_), .B2(new_n572_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n573_), .A2(new_n575_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT81), .ZN(new_n582_));
  XOR2_X1   g381(.A(G169gat), .B(G197gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n584_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT82), .Z(new_n588_));
  AND2_X1   g387(.A1(new_n562_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n576_), .A2(new_n246_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT76), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT78), .ZN(new_n593_));
  INV_X1    g392(.A(new_n246_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(new_n572_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(KEYINPUT77), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT34), .Z(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT75), .B(KEYINPUT35), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n600_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n592_), .A2(new_n595_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n603_), .A2(new_n598_), .B1(KEYINPUT36), .B2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n601_), .A2(new_n611_), .A3(new_n602_), .A4(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT37), .B1(new_n610_), .B2(new_n612_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n569_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n247_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n620_), .A2(KEYINPUT17), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(KEYINPUT79), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(KEYINPUT17), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(new_n627_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT80), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n617_), .A2(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n295_), .A2(new_n589_), .A3(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n564_), .A3(new_n549_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n587_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT109), .B1(new_n293_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT109), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n637_), .B(new_n587_), .C1(new_n288_), .C2(new_n292_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n630_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n636_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n562_), .A2(new_n613_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(new_n549_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n634_), .B1(new_n564_), .B2(new_n642_), .ZN(new_n643_));
  MUX2_X1   g442(.A(new_n634_), .B(new_n643_), .S(KEYINPUT38), .Z(G1324gat));
  NAND3_X1  g443(.A1(new_n633_), .A2(new_n565_), .A3(new_n394_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n394_), .A3(new_n641_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(new_n647_), .A3(G8gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n646_), .B2(G8gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n633_), .A2(new_n652_), .A3(new_n547_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n640_), .A2(new_n547_), .A3(new_n641_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n654_), .B2(G15gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(G22gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n633_), .A2(new_n658_), .A3(new_n554_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n640_), .A2(new_n554_), .A3(new_n641_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G22gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G22gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(new_n293_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n613_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n631_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n589_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n549_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n631_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n636_), .A2(new_n638_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n562_), .A2(new_n674_), .A3(new_n617_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n562_), .B2(new_n617_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n673_), .B(KEYINPUT44), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n549_), .A2(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n671_), .B1(new_n681_), .B2(new_n682_), .ZN(G1328gat));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n394_), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n552_), .A2(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n589_), .A2(new_n668_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n685_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT46), .B1(new_n691_), .B2(KEYINPUT110), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(new_n684_), .B2(G36gat), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n693_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n692_), .A2(new_n696_), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n679_), .A2(G43gat), .A3(new_n547_), .A4(new_n680_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n669_), .A2(new_n557_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(G43gat), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g500(.A1(new_n681_), .A2(new_n554_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G50gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n525_), .A2(G50gat), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT111), .Z(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n669_), .B2(new_n705_), .ZN(G1331gat));
  NAND4_X1  g505(.A1(new_n562_), .A2(new_n587_), .A3(new_n665_), .A4(new_n632_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n708_), .A2(KEYINPUT112), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(KEYINPUT112), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n549_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n631_), .A2(new_n588_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n641_), .A2(new_n294_), .A3(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n550_), .A2(new_n712_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n711_), .A2(new_n712_), .B1(new_n714_), .B2(new_n715_), .ZN(G1332gat));
  OR3_X1    g515(.A1(new_n707_), .A2(G64gat), .A3(new_n552_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n714_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G64gat), .B1(new_n718_), .B2(new_n552_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT48), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT48), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1333gat));
  OR3_X1    g521(.A1(new_n707_), .A2(G71gat), .A3(new_n557_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n714_), .A2(new_n547_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT49), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(new_n725_), .A3(G71gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n724_), .B2(G71gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(G1334gat));
  OR3_X1    g529(.A1(new_n707_), .A2(G78gat), .A3(new_n525_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n714_), .A2(new_n554_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(G78gat), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G78gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n293_), .A2(new_n635_), .A3(new_n672_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742_), .B2(new_n550_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n562_), .A2(new_n587_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n295_), .A2(new_n744_), .A3(new_n667_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n219_), .A3(new_n549_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1336gat));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n220_), .A3(new_n394_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n552_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n220_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT116), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n748_), .C1(new_n749_), .C2(new_n220_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n745_), .A2(new_n230_), .A3(new_n547_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n557_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n756_));
  INV_X1    g555(.A(G99gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT51), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n755_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1338gat));
  OAI211_X1 g561(.A(new_n737_), .B(new_n554_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT117), .B1(new_n763_), .B2(G106gat), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n525_), .A2(G106gat), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n764_), .A2(new_n765_), .B1(new_n745_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(G106gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT52), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n768_), .A2(new_n769_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n767_), .B(new_n775_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  NOR4_X1   g576(.A1(new_n615_), .A2(new_n616_), .A3(new_n588_), .A4(new_n631_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n291_), .A2(new_n285_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n779_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n266_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n251_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n268_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n267_), .A2(new_n785_), .A3(new_n272_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n278_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n278_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n282_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n584_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n574_), .B1(new_n578_), .B2(new_n572_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n577_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n586_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n795_), .A2(new_n587_), .B1(new_n289_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n613_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(KEYINPUT57), .A3(new_n613_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n795_), .B2(new_n801_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n794_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n282_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT58), .A3(new_n800_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n812_), .A3(new_n617_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n805_), .A2(new_n806_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n784_), .B1(new_n814_), .B2(new_n631_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n547_), .B(new_n549_), .C1(new_n553_), .C2(new_n555_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT59), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n816_), .B(new_n819_), .C1(new_n818_), .C2(new_n817_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n813_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n813_), .A2(new_n821_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n639_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n784_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n817_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n820_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n588_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G113gat), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n827_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n587_), .A2(G113gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(G1340gat));
  OAI21_X1  g633(.A(G120gat), .B1(new_n829_), .B2(new_n295_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836_));
  AOI21_X1  g635(.A(G120gat), .B1(new_n665_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT120), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n836_), .B2(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n835_), .B1(new_n832_), .B2(new_n841_), .ZN(G1341gat));
  OAI21_X1  g641(.A(G127gat), .B1(new_n829_), .B2(new_n639_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n631_), .A2(G127gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n832_), .B2(new_n844_), .ZN(G1342gat));
  INV_X1    g644(.A(new_n617_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G134gat), .B1(new_n829_), .B2(new_n846_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n613_), .A2(G134gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n832_), .B2(new_n848_), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n825_), .A2(new_n826_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n557_), .A2(new_n549_), .A3(new_n552_), .A4(new_n554_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT121), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n587_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n295_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g656(.A1(new_n853_), .A2(new_n631_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT61), .B(G155gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  INV_X1    g659(.A(G162gat), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n853_), .A2(new_n861_), .A3(new_n846_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n853_), .B2(new_n613_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n863_), .A2(KEYINPUT122), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(KEYINPUT122), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n557_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT123), .Z(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n554_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n816_), .A2(new_n867_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n870_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT125), .B1(new_n815_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n328_), .A3(new_n635_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n815_), .A2(new_n872_), .A3(new_n587_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n316_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n875_), .B1(new_n881_), .B2(new_n882_), .ZN(G1348gat));
  AOI21_X1  g682(.A(G176gat), .B1(new_n874_), .B2(new_n665_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n554_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n295_), .A2(new_n317_), .A3(new_n869_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  NOR2_X1   g686(.A1(new_n639_), .A2(new_n312_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n869_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(new_n672_), .A3(new_n889_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n874_), .A2(new_n888_), .B1(new_n890_), .B2(new_n321_), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n874_), .A2(new_n666_), .A3(new_n313_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n874_), .A2(new_n617_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(G190gat), .ZN(new_n895_));
  AOI211_X1 g694(.A(KEYINPUT126), .B(new_n322_), .C1(new_n874_), .C2(new_n617_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n892_), .B1(new_n895_), .B2(new_n896_), .ZN(G1351gat));
  NOR3_X1   g696(.A1(new_n547_), .A2(new_n552_), .A3(new_n483_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n850_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n635_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n294_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n630_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT63), .B(G211gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n899_), .B2(new_n666_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n617_), .A2(G218gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT127), .Z(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n899_), .B2(new_n911_), .ZN(G1355gat));
endmodule


