//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G43gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  INV_X1    g006(.A(KEYINPUT79), .ZN(new_n208_));
  INV_X1    g007(.A(G169gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(KEYINPUT22), .ZN(new_n210_));
  AOI21_X1  g009(.A(G176gat), .B1(new_n209_), .B2(KEYINPUT22), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT80), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n214_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT81), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(KEYINPUT81), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n221_), .A2(new_n223_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT76), .ZN(new_n235_));
  INV_X1    g034(.A(G176gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n209_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n239_), .A2(KEYINPUT78), .A3(KEYINPUT24), .A4(new_n219_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT78), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n217_), .A2(new_n218_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(KEYINPUT24), .A3(new_n238_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT24), .B1(new_n237_), .B2(new_n238_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n226_), .A2(new_n227_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OR3_X1    g046(.A1(new_n229_), .A2(KEYINPUT75), .A3(KEYINPUT26), .ZN(new_n248_));
  OR2_X1    g047(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT26), .B1(new_n229_), .B2(KEYINPUT75), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n240_), .A2(new_n244_), .A3(new_n247_), .A4(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n234_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G71gat), .B(G99gat), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n234_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n207_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n205_), .B(new_n206_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n259_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n234_), .B2(new_n254_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT83), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT31), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n260_), .A2(new_n264_), .A3(KEYINPUT83), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n267_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n265_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G64gat), .B(G92gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291_));
  INV_X1    g090(.A(G197gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(G204gat), .ZN(new_n293_));
  INV_X1    g092(.A(G204gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT85), .B1(new_n294_), .B2(G197gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(G197gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(G211gat), .A2(G218gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G211gat), .A2(G218gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n297_), .A2(new_n301_), .A3(KEYINPUT21), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT86), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT21), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(new_n293_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n292_), .A2(G204gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT21), .B1(new_n296_), .B2(new_n307_), .ZN(new_n308_));
  AND4_X1   g107(.A1(new_n304_), .A2(new_n306_), .A3(new_n300_), .A4(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n292_), .A2(G204gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n294_), .A2(G197gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n312_), .A2(KEYINPUT21), .B1(new_n298_), .B2(new_n299_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n304_), .B1(new_n313_), .B2(new_n306_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n303_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n290_), .B1(new_n255_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n306_), .A2(new_n300_), .A3(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT86), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n313_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n302_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n249_), .A2(new_n250_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n323_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n239_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n212_), .A2(G169gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n209_), .A2(KEYINPUT22), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT90), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT90), .B1(new_n326_), .B2(new_n327_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n236_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n231_), .A2(new_n219_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n324_), .A2(new_n325_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n320_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n289_), .B1(new_n316_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(new_n319_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n335_), .A2(new_n234_), .A3(new_n303_), .A4(new_n254_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n323_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n325_), .A2(new_n247_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n330_), .A2(new_n331_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n315_), .A2(new_n340_), .ZN(new_n341_));
  AND4_X1   g140(.A1(KEYINPUT20), .A2(new_n336_), .A3(new_n341_), .A4(new_n289_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n286_), .B1(new_n334_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n255_), .A2(new_n315_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(KEYINPUT20), .A3(new_n333_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n289_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n286_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n336_), .A2(new_n341_), .A3(KEYINPUT20), .A4(new_n289_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n343_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353_));
  OAI211_X1 g152(.A(KEYINPUT92), .B(new_n286_), .C1(new_n334_), .C2(new_n342_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT97), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n343_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT97), .B(new_n286_), .C1(new_n334_), .C2(new_n342_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n336_), .A2(new_n341_), .A3(KEYINPUT20), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(new_n289_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT87), .B1(new_n335_), .B2(new_n303_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n363_));
  AOI211_X1 g162(.A(new_n363_), .B(new_n302_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n332_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n255_), .B2(new_n315_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n346_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT96), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n361_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n315_), .A2(new_n363_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n335_), .A2(KEYINPUT87), .A3(new_n303_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n340_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n366_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n344_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n289_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT96), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n286_), .B1(new_n370_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n355_), .B1(new_n359_), .B2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G22gat), .B(G50gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT28), .ZN(new_n381_));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385_));
  INV_X1    g184(.A(G141gat), .ZN(new_n386_));
  INV_X1    g185(.A(G148gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT2), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n388_), .A2(new_n391_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(KEYINPUT1), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT1), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G155gat), .A3(G162gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n401_), .A3(new_n395_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n386_), .A2(new_n387_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n389_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT84), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n371_), .A2(new_n409_), .A3(new_n372_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n408_), .B1(new_n320_), .B2(new_n406_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n412_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT88), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n420_), .B2(new_n413_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n384_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n416_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n383_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n405_), .A2(new_n274_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n398_), .A2(new_n404_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT4), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n405_), .A2(new_n274_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n427_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G1gat), .B(G29gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G57gat), .B(G85gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n427_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n440_));
  OR3_X1    g239(.A1(new_n433_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n438_), .B1(new_n433_), .B2(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n379_), .A2(new_n426_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n286_), .A2(KEYINPUT32), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n334_), .B2(new_n342_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n443_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n360_), .A2(new_n289_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n369_), .B(new_n289_), .C1(new_n373_), .C2(new_n375_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n377_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n445_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n447_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n352_), .A2(new_n354_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n430_), .A2(new_n432_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n439_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n440_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(KEYINPUT94), .A3(KEYINPUT33), .A4(new_n438_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n430_), .A2(new_n427_), .A3(new_n432_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n428_), .A2(new_n429_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n438_), .B1(new_n462_), .B2(new_n439_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n442_), .A2(new_n460_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT94), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n442_), .B2(new_n460_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n454_), .A2(new_n459_), .A3(new_n467_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n453_), .A2(new_n468_), .B1(new_n425_), .B2(new_n422_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n281_), .B1(new_n444_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n443_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n423_), .A2(new_n424_), .A3(new_n383_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n383_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n280_), .B(new_n471_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(new_n379_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478_));
  INV_X1    g277(.A(G1gat), .ZN(new_n479_));
  INV_X1    g278(.A(G8gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G29gat), .B(G36gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n486_), .B(new_n489_), .Z(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(G229gat), .A3(G233gat), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n489_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n489_), .B(KEYINPUT15), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n486_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G169gat), .B(G197gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT74), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n491_), .A2(new_n496_), .A3(new_n501_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n477_), .A2(KEYINPUT98), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT98), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n464_), .A2(new_n466_), .A3(new_n459_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n354_), .B2(new_n352_), .ZN(new_n509_));
  OAI22_X1  g308(.A1(new_n509_), .A2(new_n452_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n449_), .A2(new_n448_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n365_), .A2(new_n367_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n369_), .B1(new_n512_), .B2(new_n289_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n348_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n353_), .B1(new_n343_), .B2(new_n356_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n358_), .A3(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n516_), .A2(new_n425_), .A3(new_n422_), .A4(new_n355_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n510_), .B1(new_n517_), .B2(new_n443_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n475_), .B1(new_n518_), .B2(new_n281_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n505_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n507_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n506_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G120gat), .B(G148gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT69), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT68), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G176gat), .B(G204gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT5), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT70), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n531_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G85gat), .ZN(new_n535_));
  INV_X1    g334(.A(G92gat), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n535_), .A2(new_n536_), .A3(KEYINPUT9), .ZN(new_n537_));
  XOR2_X1   g336(.A(G85gat), .B(G92gat), .Z(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(KEYINPUT9), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT10), .B(G99gat), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n534_), .B(new_n539_), .C1(G106gat), .C2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT8), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n532_), .A2(KEYINPUT67), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(G99gat), .A3(G106gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n549_), .A2(KEYINPUT66), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(KEYINPUT66), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n543_), .B(new_n545_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(G99gat), .ZN(new_n553_));
  INV_X1    g352(.A(G106gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT65), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n553_), .B(new_n554_), .C1(new_n555_), .C2(KEYINPUT7), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n557_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n548_), .A2(new_n552_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n542_), .B1(new_n560_), .B2(new_n538_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n538_), .A2(new_n542_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n534_), .B2(new_n559_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n541_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT11), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(KEYINPUT11), .ZN(new_n567_));
  XOR2_X1   g366(.A(G71gat), .B(G78gat), .Z(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n564_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n571_), .B(new_n541_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n573_), .A2(KEYINPUT12), .A3(new_n574_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT12), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n564_), .A2(new_n580_), .A3(new_n572_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n530_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n575_), .A2(new_n576_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n576_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n529_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT13), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n583_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT71), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(KEYINPUT71), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n522_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n564_), .A2(new_n493_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n489_), .B(new_n541_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n606_), .A2(new_n614_), .A3(new_n607_), .A4(new_n610_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT72), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n605_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n602_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(KEYINPUT36), .A3(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n613_), .A2(KEYINPUT72), .A3(new_n604_), .A4(new_n615_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT37), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n486_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(new_n571_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(G211gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT16), .B(G183gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT17), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n630_), .A2(KEYINPUT17), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n626_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n623_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT73), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n599_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n479_), .A3(new_n443_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n640_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n519_), .A2(new_n635_), .A3(new_n622_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n598_), .A3(new_n505_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n471_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(new_n642_), .A3(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n379_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G8gat), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT39), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n638_), .A2(new_n480_), .A3(new_n379_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n651_), .B(new_n653_), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n644_), .B2(new_n281_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT41), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n638_), .A2(new_n203_), .A3(new_n280_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n644_), .B2(new_n426_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n426_), .A2(G22gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT101), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n638_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(new_n622_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n635_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n522_), .A2(new_n598_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n443_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n598_), .A2(new_n635_), .A3(new_n505_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n477_), .B2(new_n623_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n472_), .A2(new_n473_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(new_n471_), .A3(new_n355_), .A4(new_n516_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n280_), .B1(new_n675_), .B2(new_n510_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n672_), .B(new_n623_), .C1(new_n676_), .C2(new_n475_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n671_), .B1(new_n673_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(G29gat), .A3(new_n443_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT37), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n622_), .B(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n519_), .B2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n670_), .B1(new_n685_), .B2(new_n677_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT44), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n669_), .B1(new_n682_), .B2(new_n687_), .ZN(G1328gat));
  NOR2_X1   g487(.A1(new_n647_), .A2(G36gat), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n522_), .A2(new_n598_), .A3(new_n667_), .A4(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n681_), .A2(new_n379_), .A3(new_n687_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G36gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n379_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n696_));
  AOI211_X1 g495(.A(new_n680_), .B(new_n670_), .C1(new_n685_), .C2(new_n677_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n693_), .B(G36gat), .C1(new_n696_), .C2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT46), .B(new_n692_), .C1(new_n695_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  AOI21_X1  g503(.A(G43gat), .B1(new_n668_), .B2(new_n280_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n681_), .A2(G43gat), .A3(new_n280_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n687_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n668_), .B2(new_n674_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n681_), .A2(G50gat), .A3(new_n674_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n687_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT105), .ZN(G1331gat));
  NAND3_X1  g512(.A1(new_n477_), .A2(KEYINPUT106), .A3(new_n520_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n715_), .B1(new_n519_), .B2(new_n505_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(new_n597_), .A3(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n637_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n443_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n505_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n643_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT107), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n443_), .A2(G57gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n379_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT108), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n718_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n722_), .A2(new_n379_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G64gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT48), .B(new_n725_), .C1(new_n722_), .C2(new_n379_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1333gat));
  INV_X1    g532(.A(G71gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n734_), .A3(new_n280_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n722_), .A2(new_n280_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G71gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT49), .B(new_n734_), .C1(new_n722_), .C2(new_n280_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n718_), .A2(new_n741_), .A3(new_n674_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n722_), .A2(new_n674_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(G78gat), .ZN(new_n745_));
  AOI211_X1 g544(.A(KEYINPUT50), .B(new_n741_), .C1(new_n722_), .C2(new_n674_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1335gat));
  NAND4_X1  g546(.A1(new_n714_), .A2(new_n716_), .A3(new_n597_), .A4(new_n667_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n443_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n720_), .A2(new_n635_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n685_), .B2(new_n677_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n753_), .A2(new_n535_), .A3(new_n471_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n750_), .A2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n749_), .B2(new_n379_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n753_), .A2(new_n536_), .A3(new_n647_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1337gat));
  AOI21_X1  g557(.A(new_n553_), .B1(new_n752_), .B2(new_n280_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT109), .Z(new_n760_));
  OR3_X1    g559(.A1(new_n748_), .A2(new_n540_), .A3(new_n281_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1338gat));
  NAND2_X1  g564(.A1(new_n674_), .A2(new_n554_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n748_), .A2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT111), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n554_), .B1(new_n752_), .B2(new_n674_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(KEYINPUT112), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n770_), .B2(new_n769_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT112), .B1(new_n769_), .B2(new_n770_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT53), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n768_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1339gat));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n635_), .A2(new_n505_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n583_), .A2(new_n591_), .A3(new_n588_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n591_), .B1(new_n583_), .B2(new_n588_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n593_), .A2(KEYINPUT113), .A3(new_n781_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n780_), .B1(new_n788_), .B2(new_n684_), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT54), .B(new_n623_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n578_), .A2(KEYINPUT114), .ZN(new_n794_));
  OAI22_X1  g593(.A1(KEYINPUT55), .A2(new_n582_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n793_), .A2(new_n794_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n530_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n530_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n798_), .A2(new_n588_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n501_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n494_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n495_), .B2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(new_n504_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n801_), .A2(new_n802_), .A3(KEYINPUT58), .A4(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n798_), .A2(new_n588_), .A3(new_n806_), .A4(new_n800_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n684_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT115), .B1(new_n808_), .B2(new_n809_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n798_), .A2(new_n588_), .A3(new_n505_), .A4(new_n800_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n589_), .A2(new_n806_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n665_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(KEYINPUT57), .A3(new_n665_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n812_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n791_), .B1(new_n635_), .B2(new_n820_), .ZN(new_n821_));
  NOR4_X1   g620(.A1(new_n674_), .A2(new_n379_), .A3(new_n281_), .A4(new_n471_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT59), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n815_), .B2(new_n665_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n817_), .B(new_n622_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n666_), .B1(new_n828_), .B2(new_n812_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n825_), .B(new_n822_), .C1(new_n829_), .C2(new_n791_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n824_), .A2(new_n505_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G113gat), .ZN(new_n832_));
  NOR4_X1   g631(.A1(new_n821_), .A2(G113gat), .A3(new_n520_), .A4(new_n823_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n779_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT116), .B(new_n833_), .C1(new_n831_), .C2(G113gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1340gat));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n824_), .A2(new_n597_), .A3(new_n830_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n840_), .B2(new_n839_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n820_), .A2(new_n635_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n791_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n822_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n838_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n847_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n842_), .A2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g649(.A(G127gat), .B1(new_n847_), .B2(new_n666_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n824_), .A2(new_n830_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n666_), .A2(G127gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n846_), .B2(new_n665_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n856_), .A2(KEYINPUT118), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n852_), .A2(G134gat), .A3(new_n623_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(KEYINPUT118), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(G1343gat));
  NOR3_X1   g659(.A1(new_n517_), .A2(new_n471_), .A3(new_n280_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n845_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n520_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n386_), .ZN(G1344gat));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n598_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n387_), .ZN(G1345gat));
  NOR2_X1   g665(.A1(new_n862_), .A2(new_n635_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT61), .B(G155gat), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  NOR2_X1   g668(.A1(new_n862_), .A2(new_n665_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n623_), .A2(G162gat), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n870_), .A2(G162gat), .B1(new_n862_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1347gat));
  INV_X1    g673(.A(new_n474_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n379_), .B(new_n875_), .C1(new_n829_), .C2(new_n791_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n209_), .B1(new_n877_), .B2(new_n505_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n878_), .A2(new_n879_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n505_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT120), .Z(new_n884_));
  OAI22_X1  g683(.A1(new_n881_), .A2(new_n882_), .B1(new_n876_), .B2(new_n884_), .ZN(G1348gat));
  NOR2_X1   g684(.A1(new_n876_), .A2(new_n598_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n236_), .ZN(G1349gat));
  OAI21_X1  g686(.A(new_n228_), .B1(new_n876_), .B2(new_n635_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n647_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n251_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n889_), .A2(new_n666_), .A3(new_n890_), .A4(new_n875_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n891_), .A3(KEYINPUT121), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n877_), .A2(new_n894_), .A3(new_n666_), .A4(new_n890_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n892_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n892_), .B2(new_n895_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n876_), .B2(new_n684_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n321_), .A2(new_n322_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n622_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n876_), .B2(new_n901_), .ZN(G1351gat));
  NOR3_X1   g701(.A1(new_n426_), .A2(new_n443_), .A3(new_n280_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n889_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(G197gat), .A3(new_n505_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n292_), .B1(new_n904_), .B2(new_n520_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1352gat));
  NOR2_X1   g710(.A1(new_n904_), .A2(new_n598_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT124), .B(G204gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1353gat));
  AOI21_X1  g713(.A(new_n635_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n905_), .A2(new_n915_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT125), .B(KEYINPUT126), .Z(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n916_), .B(new_n919_), .Z(G1354gat));
  XNOR2_X1  g719(.A(KEYINPUT127), .B(G218gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n904_), .A2(new_n684_), .A3(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n905_), .A2(new_n622_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n921_), .ZN(G1355gat));
endmodule


