//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_;
  XOR2_X1   g000(.A(KEYINPUT86), .B(G176gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n203_), .B1(new_n204_), .B2(KEYINPUT22), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G169gat), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n202_), .B(new_n205_), .C1(new_n203_), .C2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  MUX2_X1   g010(.A(new_n209_), .B(new_n210_), .S(new_n211_), .Z(new_n212_));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n207_), .B(new_n208_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n211_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(KEYINPUT23), .B2(new_n211_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n208_), .A2(KEYINPUT24), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  MUX2_X1   g017(.A(new_n217_), .B(KEYINPUT24), .S(new_n218_), .Z(new_n219_));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT83), .B1(new_n220_), .B2(G190gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n221_), .B(new_n222_), .C1(new_n223_), .C2(KEYINPUT83), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n216_), .A2(new_n219_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n214_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT30), .ZN(new_n227_));
  XOR2_X1   g026(.A(G15gat), .B(G43gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G227gat), .A2(G233gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT87), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n229_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT88), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT31), .Z(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G99gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT20), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT95), .B1(new_n245_), .B2(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT95), .ZN(new_n247_));
  INV_X1    g046(.A(G204gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(G197gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(G204gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT21), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT96), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(G197gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n250_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT97), .ZN(new_n258_));
  XOR2_X1   g057(.A(G211gat), .B(G218gat), .Z(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n255_), .A2(new_n250_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(KEYINPUT21), .A3(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n212_), .B1(new_n223_), .B2(new_n222_), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n208_), .B(KEYINPUT99), .Z(new_n266_));
  INV_X1    g065(.A(new_n213_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n216_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n206_), .B(KEYINPUT100), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n202_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n265_), .A2(new_n219_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n244_), .B1(new_n264_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT19), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n261_), .A2(new_n263_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n276_), .A2(KEYINPUT101), .A3(new_n226_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT101), .B1(new_n276_), .B2(new_n226_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n272_), .B(new_n275_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT20), .B1(new_n264_), .B2(new_n271_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n276_), .A2(new_n226_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n274_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT103), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n285_), .B(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n280_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n272_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n274_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n288_), .B(KEYINPUT107), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(KEYINPUT27), .B(new_n289_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296_));
  INV_X1    g095(.A(new_n289_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n288_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT108), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n295_), .A2(new_n299_), .A3(KEYINPUT108), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(KEYINPUT89), .A2(G155gat), .A3(G162gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(G155gat), .B2(G162gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT92), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n309_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT91), .ZN(new_n313_));
  OR2_X1    g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n314_), .A2(KEYINPUT3), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n313_), .B(new_n317_), .C1(KEYINPUT3), .C2(new_n314_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n310_), .A2(new_n311_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n307_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(KEYINPUT1), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(KEYINPUT1), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT90), .Z(new_n324_));
  OAI211_X1 g123(.A(new_n316_), .B(new_n314_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT94), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n276_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT98), .ZN(new_n331_));
  INV_X1    g130(.A(G228gat), .ZN(new_n332_));
  INV_X1    g131(.A(G233gat), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n331_), .B(new_n336_), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n329_), .B(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n339_));
  XOR2_X1   g138(.A(G22gat), .B(G50gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT28), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n339_), .B(new_n341_), .Z(new_n342_));
  OR2_X1    g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n342_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n302_), .A2(new_n303_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n243_), .B1(new_n347_), .B2(KEYINPUT109), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT109), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n302_), .A2(new_n303_), .A3(new_n349_), .A4(new_n346_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n242_), .A2(new_n346_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n300_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n348_), .A2(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n319_), .A2(new_n235_), .A3(new_n325_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n236_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n326_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT105), .Z(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT104), .B(KEYINPUT4), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n326_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n356_), .B2(KEYINPUT4), .ZN(new_n362_));
  INV_X1    g161(.A(new_n357_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT0), .ZN(new_n367_));
  INV_X1    g166(.A(G57gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n359_), .A2(new_n364_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n353_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n242_), .A2(new_n345_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT33), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n362_), .A2(new_n357_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n356_), .A2(new_n363_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n371_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n297_), .A2(new_n298_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT106), .B1(new_n374_), .B2(new_n379_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n374_), .A2(KEYINPUT106), .A3(new_n379_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n385_), .B(new_n386_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n288_), .A2(KEYINPUT32), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n279_), .A2(new_n282_), .A3(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n375_), .B(new_n391_), .C1(new_n292_), .C2(new_n390_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n378_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n376_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT71), .ZN(new_n395_));
  XOR2_X1   g194(.A(G71gat), .B(G78gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(G57gat), .B(G64gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n396_), .B1(KEYINPUT11), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(KEYINPUT11), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G57gat), .B(G64gat), .Z(new_n402_));
  INV_X1    g201(.A(KEYINPUT11), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n402_), .A2(new_n396_), .A3(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT12), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT9), .ZN(new_n408_));
  INV_X1    g207(.A(G92gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n370_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G85gat), .A2(G92gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n408_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT65), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(G85gat), .A2(G92gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G85gat), .A2(G92gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT9), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT65), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n413_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT67), .ZN(new_n422_));
  OR2_X1    g221(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n423_));
  OR2_X1    g222(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT66), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G99gat), .A2(G106gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n434_));
  NAND3_X1  g233(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n427_), .A2(new_n430_), .A3(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n421_), .A2(new_n422_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n422_), .B1(new_n421_), .B2(new_n437_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n416_), .A2(new_n417_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT8), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n430_), .A2(new_n436_), .ZN(new_n444_));
  INV_X1    g243(.A(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(G106gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(KEYINPUT68), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT7), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(new_n445_), .A3(new_n446_), .A4(KEYINPUT68), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n443_), .B1(new_n444_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT68), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(G99gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n449_), .B1(new_n455_), .B2(new_n446_), .ZN(new_n456_));
  NOR4_X1   g255(.A1(new_n454_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT69), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n433_), .A2(new_n435_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n448_), .A2(new_n461_), .A3(new_n450_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n441_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n453_), .B1(new_n464_), .B2(KEYINPUT8), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n407_), .B1(new_n440_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n404_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n402_), .A2(new_n403_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n399_), .A3(new_n396_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n471_), .A3(KEYINPUT70), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n412_), .A2(new_n414_), .A3(KEYINPUT65), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n419_), .B1(new_n418_), .B2(new_n413_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n444_), .A2(new_n427_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT67), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n421_), .A2(new_n422_), .A3(new_n437_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n430_), .A2(new_n436_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n442_), .B(new_n441_), .C1(new_n481_), .C2(new_n451_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n441_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n459_), .B1(new_n451_), .B2(KEYINPUT69), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n462_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n482_), .B1(new_n485_), .B2(new_n442_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n473_), .B1(new_n480_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n466_), .B1(new_n487_), .B2(KEYINPUT12), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n486_), .A3(new_n473_), .ZN(new_n489_));
  INV_X1    g288(.A(G230gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(new_n333_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n395_), .B1(new_n488_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n468_), .A2(new_n472_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n440_), .B2(new_n465_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT12), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n464_), .A2(KEYINPUT8), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n499_), .A2(new_n482_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n491_), .B1(new_n500_), .B2(new_n473_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n498_), .A2(new_n501_), .A3(KEYINPUT71), .A4(new_n466_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n494_), .A2(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n480_), .A2(new_n486_), .A3(new_n473_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n491_), .B1(new_n504_), .B2(new_n487_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(KEYINPUT72), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G120gat), .B(G148gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(new_n248_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT5), .B(G176gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n494_), .A2(new_n505_), .A3(new_n502_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n506_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n503_), .A2(new_n516_), .A3(new_n505_), .A4(new_n510_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT73), .B1(new_n512_), .B2(new_n511_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n515_), .A2(new_n519_), .A3(KEYINPUT13), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G113gat), .B(G141gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G169gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(new_n245_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528_));
  INV_X1    g327(.A(G1gat), .ZN(new_n529_));
  INV_X1    g328(.A(G8gat), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT14), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT79), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT79), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n534_), .A3(new_n531_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G1gat), .B(G8gat), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G36gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(G43gat), .B(G50gat), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT74), .ZN(new_n545_));
  INV_X1    g344(.A(G29gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G43gat), .B(G50gat), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n546_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n543_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n549_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n547_), .A2(new_n548_), .ZN(new_n555_));
  OAI21_X1  g354(.A(G29gat), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(G36gat), .A3(new_n550_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n553_), .A2(KEYINPUT15), .A3(new_n557_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n542_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n551_), .A2(new_n552_), .A3(new_n543_), .ZN(new_n563_));
  AOI21_X1  g362(.A(G36gat), .B1(new_n556_), .B2(new_n550_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n542_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n562_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n567_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n558_), .A2(new_n541_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n553_), .A2(new_n557_), .B1(new_n540_), .B2(new_n539_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n527_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n573_), .B(new_n527_), .C1(new_n562_), .C2(new_n568_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n524_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n560_), .A2(new_n561_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n442_), .B1(new_n463_), .B2(new_n441_), .ZN(new_n581_));
  OAI22_X1  g380(.A1(new_n581_), .A2(new_n453_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n500_), .A2(new_n565_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n583_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n586_), .A2(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n583_), .A2(new_n593_), .A3(new_n588_), .A4(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT78), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(KEYINPUT78), .A3(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT36), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n592_), .A2(new_n594_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(new_n604_), .A3(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n602_), .B(KEYINPUT76), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT37), .B1(new_n607_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT77), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT77), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n614_), .B(KEYINPUT37), .C1(new_n607_), .C2(new_n611_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n609_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n541_), .B(new_n617_), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n473_), .ZN(new_n619_));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT17), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n619_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n405_), .B(KEYINPUT80), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n618_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n624_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n618_), .A2(new_n627_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n616_), .A2(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n394_), .A2(new_n579_), .A3(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n529_), .A3(new_n375_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT38), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n603_), .A2(new_n608_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n394_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n633_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n579_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n375_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n637_), .A2(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n389_), .A2(new_n392_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n648_), .A2(new_n378_), .B1(new_n353_), .B2(new_n375_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n302_), .A2(new_n303_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n638_), .A4(new_n642_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n647_), .B1(new_n651_), .B2(G8gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n647_), .A3(G8gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n635_), .A2(new_n530_), .A3(new_n650_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT110), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n659_));
  INV_X1    g458(.A(new_n654_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n659_), .B(new_n656_), .C1(new_n660_), .C2(new_n652_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(KEYINPUT40), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n659_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n661_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(G1325gat));
  INV_X1    g466(.A(G15gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n635_), .A2(new_n668_), .A3(new_n242_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G15gat), .B1(new_n643_), .B2(new_n243_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n635_), .A2(new_n675_), .A3(new_n345_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G22gat), .B1(new_n643_), .B2(new_n346_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT111), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT111), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n679_), .B(G22gat), .C1(new_n643_), .C2(new_n346_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n678_), .A2(KEYINPUT42), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT42), .B1(new_n678_), .B2(new_n680_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n681_), .B2(new_n682_), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n394_), .A2(new_n638_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n579_), .A2(new_n633_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n375_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n609_), .A2(new_n615_), .A3(new_n613_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n689_), .B(new_n690_), .C1(new_n376_), .C2(new_n393_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(new_n649_), .B2(new_n690_), .ZN(new_n693_));
  OAI211_X1 g492(.A(KEYINPUT44), .B(new_n685_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(G29gat), .A3(new_n375_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n685_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n688_), .B1(new_n695_), .B2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  INV_X1    g499(.A(new_n650_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n685_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n394_), .B2(new_n616_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n691_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n701_), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n543_), .B1(new_n705_), .B2(new_n698_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n684_), .A2(new_n543_), .A3(new_n650_), .A4(new_n685_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n707_), .B(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n700_), .B1(new_n706_), .B2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n704_), .A2(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n694_), .A2(new_n650_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G36gat), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n707_), .B(new_n708_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(KEYINPUT46), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n716_), .ZN(G1329gat));
  INV_X1    g516(.A(G43gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n686_), .B2(new_n243_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n694_), .A2(G43gat), .A3(new_n242_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n712_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT47), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n723_), .B(new_n719_), .C1(new_n720_), .C2(new_n712_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1330gat));
  OR3_X1    g524(.A1(new_n686_), .A2(G50gat), .A3(new_n346_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n694_), .A2(new_n345_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT113), .B(G50gat), .C1(new_n712_), .C2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n698_), .A2(new_n345_), .A3(new_n694_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT113), .B1(new_n730_), .B2(G50gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n729_), .B2(new_n731_), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n524_), .A2(new_n578_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n640_), .A2(new_n633_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n644_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n733_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n394_), .A2(new_n634_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n368_), .A3(new_n375_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n740_), .A3(new_n650_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G64gat), .B1(new_n734_), .B2(new_n701_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT48), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT48), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n746_), .A3(new_n242_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G71gat), .B1(new_n734_), .B2(new_n243_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n737_), .A2(new_n752_), .A3(new_n345_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G78gat), .B1(new_n734_), .B2(new_n346_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT50), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT50), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n703_), .A2(new_n691_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n736_), .A2(new_n633_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n644_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n684_), .A2(new_n759_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n763_), .B2(new_n650_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n760_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n650_), .A2(G92gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT114), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n767_), .B2(new_n769_), .ZN(G1337gat));
  NAND3_X1  g569(.A1(new_n758_), .A2(new_n242_), .A3(new_n759_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G99gat), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n242_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n763_), .A2(new_n773_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  OR2_X1    g574(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(G1338gat));
  NAND4_X1  g576(.A1(new_n763_), .A2(new_n345_), .A3(new_n424_), .A4(new_n426_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n345_), .B(new_n759_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n778_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NAND2_X1  g586(.A1(new_n348_), .A2(new_n350_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n375_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n577_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n406_), .B1(new_n480_), .B2(new_n486_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT116), .B1(new_n795_), .B2(new_n489_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT12), .B1(new_n582_), .B2(new_n495_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NOR4_X1   g597(.A1(new_n797_), .A2(new_n504_), .A3(new_n794_), .A4(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n491_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n494_), .A2(new_n801_), .A3(new_n502_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n488_), .A2(new_n493_), .A3(new_n801_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT117), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n511_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n793_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n805_), .B2(new_n511_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n792_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n494_), .A2(new_n801_), .A3(new_n502_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n466_), .B(new_n489_), .C1(new_n487_), .C2(KEYINPUT12), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n798_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n498_), .A2(KEYINPUT116), .A3(new_n489_), .A4(new_n466_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n492_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n813_), .A2(new_n817_), .A3(new_n803_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n807_), .B1(new_n818_), .B2(new_n510_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(new_n793_), .A3(KEYINPUT118), .A4(new_n809_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n567_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n527_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n566_), .A2(new_n570_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n821_), .B(new_n822_), .C1(new_n562_), .C2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n575_), .A2(new_n824_), .A3(KEYINPUT119), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT119), .B1(new_n575_), .B2(new_n824_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n812_), .A2(new_n820_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n638_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n827_), .B1(new_n518_), .B2(new_n517_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n815_), .A2(new_n816_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n803_), .B1(new_n835_), .B2(new_n491_), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n806_), .B(new_n510_), .C1(new_n836_), .C2(new_n802_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n511_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n834_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n834_), .B(KEYINPUT58), .C1(new_n837_), .C2(new_n838_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(new_n690_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n833_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n830_), .B2(new_n638_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT121), .B1(new_n847_), .B2(new_n843_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n633_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n634_), .A2(new_n578_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n850_), .A2(new_n524_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n850_), .B2(new_n524_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n791_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n819_), .A2(new_n809_), .A3(new_n793_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n828_), .B1(new_n856_), .B2(new_n792_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n639_), .B1(new_n857_), .B2(new_n820_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n843_), .B1(new_n858_), .B2(KEYINPUT57), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n858_), .B2(KEYINPUT57), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n831_), .A2(KEYINPUT120), .A3(new_n832_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n854_), .B1(new_n863_), .B2(new_n641_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT59), .B1(new_n864_), .B2(new_n790_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n855_), .A2(new_n865_), .A3(new_n578_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G113gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n864_), .A2(new_n790_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n577_), .A2(G113gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n867_), .B1(new_n869_), .B2(new_n870_), .ZN(G1340gat));
  NOR2_X1   g670(.A1(new_n524_), .A2(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(KEYINPUT60), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n524_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n865_), .A4(new_n855_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(KEYINPUT60), .B2(new_n873_), .ZN(G1341gat));
  NAND3_X1  g676(.A1(new_n855_), .A2(new_n865_), .A3(new_n633_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G127gat), .ZN(new_n879_));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n868_), .A2(new_n880_), .A3(new_n633_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT122), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n879_), .A2(new_n884_), .A3(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1342gat));
  NAND3_X1  g685(.A1(new_n855_), .A2(new_n865_), .A3(new_n690_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G134gat), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n638_), .A2(G134gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n869_), .B2(new_n889_), .ZN(G1343gat));
  INV_X1    g689(.A(new_n864_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n701_), .A2(new_n375_), .A3(new_n351_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n578_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n874_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g697(.A1(new_n893_), .A2(new_n641_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT61), .B(G155gat), .Z(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  OAI21_X1  g700(.A(G162gat), .B1(new_n893_), .B2(new_n616_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n638_), .A2(G162gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n893_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT123), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n902_), .B(new_n906_), .C1(new_n893_), .C2(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n858_), .A2(KEYINPUT57), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n841_), .A2(new_n690_), .A3(new_n842_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n845_), .B(new_n911_), .C1(new_n858_), .C2(KEYINPUT57), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n848_), .A2(new_n910_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n854_), .B1(new_n913_), .B2(new_n641_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n701_), .A2(new_n375_), .A3(new_n243_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n346_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n914_), .A2(new_n577_), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n909_), .B1(new_n917_), .B2(new_n204_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n269_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n916_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n578_), .B(new_n920_), .C1(new_n849_), .C2(new_n854_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n918_), .A2(new_n919_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT124), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n918_), .A2(new_n919_), .A3(new_n925_), .A4(new_n922_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1348gat));
  NOR2_X1   g726(.A1(new_n914_), .A2(new_n916_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n874_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n864_), .A2(new_n345_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n915_), .A2(new_n874_), .A3(G176gat), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n929_), .A2(new_n202_), .B1(new_n930_), .B2(new_n931_), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n633_), .A3(new_n915_), .ZN(new_n933_));
  INV_X1    g732(.A(G183gat), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n641_), .A2(new_n222_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n934_), .B1(new_n928_), .B2(new_n935_), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n928_), .A2(new_n223_), .A3(new_n639_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n914_), .A2(new_n616_), .A3(new_n916_), .ZN(new_n938_));
  INV_X1    g737(.A(G190gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(G1351gat));
  NAND2_X1  g739(.A1(new_n644_), .A2(new_n351_), .ZN(new_n941_));
  XOR2_X1   g740(.A(new_n941_), .B(KEYINPUT125), .Z(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n650_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n864_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n578_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g745(.A(new_n944_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n524_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n248_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT126), .B(G204gat), .Z(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n948_), .B2(new_n951_), .ZN(G1353gat));
  XOR2_X1   g751(.A(KEYINPUT63), .B(G211gat), .Z(new_n953_));
  NOR3_X1   g752(.A1(new_n947_), .A2(new_n641_), .A3(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n944_), .B2(new_n633_), .ZN(new_n956_));
  OR3_X1    g755(.A1(new_n954_), .A2(new_n956_), .A3(KEYINPUT127), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT127), .B1(new_n954_), .B2(new_n956_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1354gat));
  OR3_X1    g758(.A1(new_n947_), .A2(G218gat), .A3(new_n638_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G218gat), .B1(new_n947_), .B2(new_n616_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1355gat));
endmodule


