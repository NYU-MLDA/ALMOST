//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT9), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n210_), .A2(KEYINPUT64), .A3(new_n219_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G29gat), .B(G36gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(KEYINPUT15), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT35), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G232gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n220_), .A2(new_n228_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n233_), .A2(new_n229_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n227_), .A2(new_n238_), .A3(new_n234_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G190gat), .B(G218gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G134gat), .B(G162gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT36), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT69), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n242_), .B(KEYINPUT36), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT70), .ZN(new_n247_));
  INV_X1    g046(.A(new_n239_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n238_), .B1(new_n227_), .B2(new_n234_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n237_), .A2(new_n251_), .A3(new_n239_), .A4(new_n243_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT37), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(KEYINPUT71), .B(new_n247_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n244_), .A4(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n254_), .A2(KEYINPUT73), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT73), .B1(new_n254_), .B2(new_n259_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G1gat), .ZN(new_n263_));
  INV_X1    g062(.A(G8gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT14), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n266_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G15gat), .B(G22gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G8gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n271_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n267_), .A2(new_n273_), .A3(new_n268_), .A4(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G231gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G57gat), .B(G64gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G71gat), .B(G78gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n279_), .A2(new_n281_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n277_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G127gat), .B(G155gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G183gat), .B(G211gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT77), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n287_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT78), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n287_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n287_), .A2(new_n298_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n292_), .B(KEYINPUT17), .Z(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n262_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G120gat), .B(G148gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(G176gat), .B(G204gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G230gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n286_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n222_), .A2(new_n223_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT65), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n222_), .A2(new_n315_), .A3(new_n223_), .A4(new_n312_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n222_), .A2(new_n223_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(new_n286_), .ZN(new_n320_));
  AOI211_X1 g119(.A(KEYINPUT66), .B(new_n312_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n311_), .B1(new_n317_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n220_), .A2(KEYINPUT12), .A3(new_n286_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n312_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n324_), .B(new_n313_), .C1(new_n325_), .C2(KEYINPUT12), .ZN(new_n326_));
  INV_X1    g125(.A(new_n311_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n310_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n223_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT64), .B1(new_n210_), .B2(new_n219_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n286_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT66), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n318_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n314_), .A4(new_n316_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n327_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n313_), .A2(new_n324_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n339_), .A3(new_n311_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n340_), .A3(new_n309_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n329_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT13), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n329_), .A2(new_n341_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT13), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n304_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT80), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT21), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  AND2_X1   g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G211gat), .B(G218gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G211gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(G218gat), .ZN(new_n359_));
  INV_X1    g158(.A(G218gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(G211gat), .ZN(new_n361_));
  OAI22_X1  g160(.A1(new_n359_), .A2(new_n361_), .B1(new_n354_), .B2(new_n353_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n351_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT21), .B1(new_n355_), .B2(new_n356_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT84), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(G183gat), .A3(G190gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT23), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(G183gat), .B2(G190gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n366_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT22), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(G169gat), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(KEYINPUT22), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT93), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G176gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(KEYINPUT22), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT93), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n374_), .A2(new_n375_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n368_), .A2(new_n370_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT23), .ZN(new_n389_));
  NOR3_X1   g188(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT24), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(G169gat), .B2(G176gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n378_), .A2(new_n381_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n367_), .A2(new_n372_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n389_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT26), .B(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n399_));
  INV_X1    g198(.A(G183gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(KEYINPUT25), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(G183gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n399_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(G183gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(KEYINPUT25), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT92), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n398_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n396_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n365_), .B1(new_n387_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n389_), .A2(new_n366_), .A3(new_n395_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n382_), .A2(new_n383_), .A3(new_n381_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT85), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n382_), .A2(new_n383_), .A3(new_n414_), .A4(new_n381_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n416_), .A3(new_n375_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT25), .B1(new_n400_), .B2(KEYINPUT83), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n397_), .B(new_n418_), .C1(KEYINPUT83), .C2(new_n405_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n394_), .C1(new_n373_), .C2(new_n371_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n417_), .B(new_n420_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n410_), .A2(new_n421_), .A3(KEYINPUT20), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n417_), .A2(new_n420_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n365_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n407_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT92), .B1(new_n405_), .B2(new_n406_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n397_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n395_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n388_), .B2(KEYINPUT23), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n433_), .A3(new_n394_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n374_), .A2(new_n386_), .A3(new_n375_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n434_), .B(new_n435_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n425_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n428_), .A2(new_n436_), .A3(KEYINPUT20), .A4(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n426_), .A2(KEYINPUT94), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT94), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n422_), .A2(new_n440_), .A3(new_n425_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G8gat), .B(G36gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT96), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n439_), .A2(new_n447_), .A3(new_n441_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n442_), .A2(KEYINPUT96), .A3(new_n448_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G127gat), .B(G134gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G113gat), .B(G120gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G141gat), .ZN(new_n460_));
  INV_X1    g259(.A(G148gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G141gat), .A2(G148gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT87), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G155gat), .A3(G162gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G155gat), .ZN(new_n470_));
  INV_X1    g269(.A(G162gat), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n469_), .A2(KEYINPUT1), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT1), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n464_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n471_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n469_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT88), .ZN(new_n479_));
  NAND3_X1  g278(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n477_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n459_), .B1(new_n475_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n478_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT2), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n463_), .A2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n490_), .B(new_n480_), .C1(new_n462_), .C2(KEYINPUT3), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n469_), .B(new_n476_), .C1(new_n488_), .C2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n469_), .A2(KEYINPUT1), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n493_), .A2(new_n476_), .A3(new_n474_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n492_), .B(new_n458_), .C1(new_n494_), .C2(new_n464_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G225gat), .A2(G233gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n486_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G29gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G85gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT0), .B(G57gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  AND3_X1   g300(.A1(new_n486_), .A2(new_n495_), .A3(KEYINPUT4), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n459_), .B(new_n503_), .C1(new_n475_), .C2(new_n485_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n496_), .B(KEYINPUT97), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n497_), .B(new_n501_), .C1(new_n502_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n486_), .A2(new_n495_), .A3(KEYINPUT4), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n501_), .B1(new_n510_), .B2(new_n497_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n508_), .A2(new_n511_), .A3(KEYINPUT99), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT99), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n497_), .B1(new_n502_), .B2(new_n506_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n501_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n513_), .B1(new_n516_), .B2(new_n507_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT29), .B1(new_n475_), .B2(new_n485_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n365_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n365_), .A3(new_n521_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G78gat), .B(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT90), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n475_), .A2(new_n485_), .A3(KEYINPUT29), .ZN(new_n529_));
  XOR2_X1   g328(.A(G22gat), .B(G50gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT28), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n529_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n524_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n527_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n535_), .A2(new_n532_), .A3(new_n527_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n449_), .A2(KEYINPUT27), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT100), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n428_), .A2(KEYINPUT20), .A3(new_n436_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n425_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n410_), .A2(new_n421_), .A3(KEYINPUT20), .A4(new_n437_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n542_), .B1(new_n546_), .B2(new_n447_), .ZN(new_n547_));
  AOI211_X1 g346(.A(KEYINPUT100), .B(new_n448_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n518_), .B(new_n540_), .C1(new_n541_), .C2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT102), .B1(new_n455_), .B2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n541_), .A2(new_n549_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n539_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n528_), .A2(new_n532_), .B1(new_n535_), .B2(new_n527_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT99), .B1(new_n508_), .B2(new_n511_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n516_), .A2(new_n513_), .A3(new_n507_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT102), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n552_), .A2(new_n553_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n509_), .A2(new_n496_), .A3(new_n504_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n486_), .A2(new_n495_), .A3(new_n505_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n515_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n507_), .A2(new_n566_), .A3(KEYINPUT33), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT33), .B1(new_n507_), .B2(new_n566_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n546_), .A2(KEYINPUT32), .A3(new_n448_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(new_n511_), .B2(new_n508_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n448_), .A2(KEYINPUT32), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n442_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n556_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n551_), .A2(new_n562_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n427_), .B(KEYINPUT30), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G227gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(G15gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(G71gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(G99gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n577_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(new_n459_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT86), .B(G43gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT31), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n576_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT103), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n589_), .A2(new_n559_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n552_), .A2(new_n553_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n540_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT103), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n576_), .A2(new_n596_), .A3(new_n589_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n275_), .B(new_n226_), .Z(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n228_), .A2(new_n275_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n272_), .A2(new_n226_), .A3(new_n274_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(new_n600_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n599_), .A2(new_n601_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G113gat), .B(G141gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT82), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G169gat), .B(G197gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT81), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n605_), .B(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n598_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n350_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n263_), .A3(new_n559_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n614_), .B1(KEYINPUT105), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n616_), .B1(new_n617_), .B2(KEYINPUT38), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n256_), .A2(new_n257_), .A3(new_n244_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n598_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n611_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n347_), .A2(new_n303_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n518_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT104), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n614_), .A2(KEYINPUT105), .A3(new_n615_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n618_), .A2(new_n625_), .A3(new_n626_), .ZN(G1324gat));
  NAND3_X1  g426(.A1(new_n613_), .A2(new_n264_), .A3(new_n593_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n620_), .A2(new_n593_), .A3(new_n622_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(G8gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(G8gat), .A3(new_n629_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n628_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n623_), .B2(new_n589_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT41), .Z(new_n638_));
  INV_X1    g437(.A(new_n589_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n613_), .A2(new_n579_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1326gat));
  OAI21_X1  g440(.A(G22gat), .B1(new_n623_), .B2(new_n556_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT42), .ZN(new_n643_));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n613_), .A2(new_n644_), .A3(new_n540_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1327gat));
  INV_X1    g445(.A(new_n303_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n347_), .A2(new_n619_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n612_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n559_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n597_), .A2(new_n595_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n596_), .B1(new_n576_), .B2(new_n589_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n262_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n262_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n343_), .A2(new_n303_), .A3(new_n611_), .A4(new_n346_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n664_), .B(new_n661_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n559_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n651_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(KEYINPUT109), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(KEYINPUT109), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT110), .Z(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n666_), .B2(new_n593_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n676_));
  INV_X1    g475(.A(new_n593_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n649_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n676_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n612_), .A2(new_n648_), .A3(new_n681_), .A4(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n671_), .B(new_n673_), .C1(new_n675_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n673_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n657_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n656_), .B1(new_n598_), .B2(new_n262_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n662_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n664_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n662_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n593_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n683_), .B1(new_n691_), .B2(G36gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n685_), .B1(new_n692_), .B2(new_n670_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n684_), .A2(new_n693_), .ZN(G1329gat));
  AOI21_X1  g493(.A(G43gat), .B1(new_n650_), .B2(new_n639_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n639_), .A2(G43gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n666_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1330gat));
  NOR3_X1   g498(.A1(new_n663_), .A2(new_n665_), .A3(new_n556_), .ZN(new_n700_));
  INV_X1    g499(.A(G50gat), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n556_), .A2(G50gat), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT112), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n700_), .A2(new_n701_), .B1(new_n649_), .B2(new_n703_), .ZN(G1331gat));
  NAND4_X1  g503(.A1(new_n620_), .A2(new_n647_), .A3(new_n621_), .A4(new_n347_), .ZN(new_n705_));
  INV_X1    g504(.A(G57gat), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n518_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n348_), .A2(new_n611_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n598_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n304_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n518_), .B1(new_n710_), .B2(KEYINPUT113), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(KEYINPUT113), .B2(new_n710_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n712_), .B2(new_n706_), .ZN(G1332gat));
  OAI21_X1  g512(.A(G64gat), .B1(new_n705_), .B2(new_n677_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT48), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n677_), .A2(G64gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n710_), .B2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n705_), .B2(new_n589_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT49), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(G71gat), .C1(new_n705_), .C2(new_n589_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  OR3_X1    g521(.A1(new_n710_), .A2(G71gat), .A3(new_n589_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(KEYINPUT114), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n705_), .B2(new_n556_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n556_), .A2(G78gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n710_), .B2(new_n731_), .ZN(G1335gat));
  NOR3_X1   g531(.A1(new_n348_), .A2(new_n647_), .A3(new_n611_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n658_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n518_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n647_), .A2(new_n619_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n709_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n211_), .A3(new_n559_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n735_), .A2(new_n739_), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n734_), .B2(new_n677_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n212_), .A3(new_n593_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  NAND2_X1  g542(.A1(new_n639_), .A2(new_n215_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n737_), .A2(new_n744_), .B1(KEYINPUT115), .B2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n658_), .A2(new_n733_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n639_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(G99gat), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n745_), .A2(KEYINPUT115), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(G1338gat));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n556_), .A2(G106gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n738_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n753_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT116), .B1(new_n737_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n216_), .B1(new_n747_), .B2(new_n540_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n734_), .A2(new_n556_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n762_), .A2(new_n216_), .A3(new_n759_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT53), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n758_), .A2(new_n760_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n759_), .B1(new_n762_), .B2(new_n216_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n765_), .A2(new_n766_), .A3(new_n767_), .A4(new_n757_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n328_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n326_), .A2(new_n770_), .A3(new_n327_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n310_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT56), .B(new_n310_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n609_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT119), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n599_), .A2(new_n600_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n609_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(KEYINPUT119), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n602_), .A2(new_n603_), .A3(new_n601_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n605_), .A2(new_n609_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n341_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT58), .B1(new_n778_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n254_), .A2(new_n259_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT73), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n254_), .A2(KEYINPUT73), .A3(new_n259_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT122), .B1(new_n790_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n311_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n340_), .B1(new_n797_), .B2(new_n770_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n773_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n310_), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n775_), .B(new_n309_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n789_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n262_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n778_), .A2(KEYINPUT58), .A3(new_n789_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n796_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n619_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n341_), .A2(new_n611_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n802_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n776_), .A2(KEYINPUT118), .A3(new_n777_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n344_), .B2(new_n788_), .ZN(new_n817_));
  AOI211_X1 g616(.A(KEYINPUT120), .B(new_n787_), .C1(new_n329_), .C2(new_n341_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n810_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n809_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(KEYINPUT57), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n303_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n348_), .A2(new_n647_), .A3(new_n795_), .A4(new_n621_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n594_), .A2(new_n639_), .A3(new_n559_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n611_), .B(new_n341_), .C1(new_n777_), .C2(KEYINPUT118), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n801_), .A2(new_n802_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(KEYINPUT118), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT120), .B1(new_n342_), .B2(new_n787_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n344_), .A2(new_n816_), .A3(new_n788_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n619_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT121), .B1(new_n820_), .B2(KEYINPUT57), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n809_), .A4(new_n821_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n827_), .B1(new_n845_), .B2(new_n303_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n831_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n833_), .B1(new_n847_), .B2(new_n830_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n621_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n303_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n828_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n832_), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n852_), .A2(G113gat), .A3(new_n621_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n848_), .B2(new_n348_), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n348_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n847_), .B(new_n857_), .C1(KEYINPUT60), .C2(new_n856_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(G1341gat));
  OAI21_X1  g658(.A(G127gat), .B1(new_n848_), .B2(new_n303_), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n852_), .A2(G127gat), .A3(new_n303_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n847_), .B2(new_n810_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n848_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT123), .B(G134gat), .Z(new_n865_));
  NOR2_X1   g664(.A1(new_n795_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n864_), .B2(new_n866_), .ZN(G1343gat));
  NOR4_X1   g666(.A1(new_n639_), .A2(new_n518_), .A3(new_n556_), .A4(new_n593_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n851_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n621_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n460_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n348_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n461_), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n869_), .A2(new_n303_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n869_), .B2(new_n795_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n810_), .A2(new_n471_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n869_), .B2(new_n878_), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n592_), .A2(new_n593_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n829_), .A2(new_n556_), .A3(new_n611_), .A4(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  AND4_X1   g683(.A1(new_n880_), .A2(new_n883_), .A3(new_n884_), .A4(G169gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n378_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n883_), .A2(new_n886_), .B1(new_n880_), .B2(new_n884_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n829_), .A2(new_n556_), .A3(new_n882_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n611_), .A2(new_n380_), .A3(new_n385_), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT125), .Z(new_n890_));
  OAI22_X1  g689(.A1(new_n885_), .A2(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(G1348gat));
  OR2_X1    g690(.A1(new_n888_), .A2(new_n348_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n846_), .A2(new_n540_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n348_), .A2(new_n381_), .A3(new_n881_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n892_), .A2(new_n381_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n881_), .A2(new_n303_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n407_), .A3(new_n404_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n540_), .B(new_n897_), .C1(new_n824_), .C2(new_n828_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n893_), .A2(new_n896_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n400_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n888_), .B2(new_n795_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n810_), .A2(new_n397_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n888_), .B2(new_n902_), .ZN(G1351gat));
  NAND3_X1  g702(.A1(new_n589_), .A2(new_n560_), .A3(new_n593_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n851_), .A2(KEYINPUT126), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n846_), .B2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G197gat), .B1(new_n909_), .B2(new_n611_), .ZN(new_n910_));
  INV_X1    g709(.A(G197gat), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n911_), .B(new_n621_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1352gat));
  AOI21_X1  g712(.A(KEYINPUT126), .B1(new_n851_), .B2(new_n905_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n846_), .A2(new_n907_), .A3(new_n904_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n347_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G204gat), .ZN(new_n917_));
  INV_X1    g716(.A(G204gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n909_), .A2(new_n918_), .A3(new_n347_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1353gat));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n647_), .B1(new_n923_), .B2(new_n358_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n922_), .B1(new_n909_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n922_), .ZN(new_n927_));
  AOI211_X1 g726(.A(new_n927_), .B(new_n924_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1354gat));
  NAND3_X1  g728(.A1(new_n909_), .A2(new_n360_), .A3(new_n810_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n795_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n360_), .B2(new_n931_), .ZN(G1355gat));
endmodule


