//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n204_));
  INV_X1    g003(.A(G22gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT76), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G15gat), .ZN(new_n207_));
  INV_X1    g006(.A(G15gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT76), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(KEYINPUT76), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(G15gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(G22gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(G1gat), .B2(G8gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n204_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  AOI211_X1 g017(.A(KEYINPUT77), .B(new_n216_), .C1(new_n210_), .C2(new_n213_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n203_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n213_), .ZN(new_n221_));
  AOI21_X1  g020(.A(G22gat), .B1(new_n211_), .B2(new_n212_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n217_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT77), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n214_), .A2(new_n204_), .A3(new_n217_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n202_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G29gat), .B(G36gat), .Z(new_n228_));
  XOR2_X1   g027(.A(G43gat), .B(G50gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT15), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT81), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236_));
  INV_X1    g035(.A(new_n230_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n227_), .B2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n220_), .A2(new_n226_), .A3(KEYINPUT79), .A4(new_n230_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n235_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n230_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n233_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n249_), .A2(KEYINPUT80), .A3(new_n233_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n241_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G169gat), .B(G197gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n241_), .B(new_n254_), .C1(new_n248_), .C2(new_n250_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G78gat), .B(G106gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT93), .Z(new_n261_));
  NAND2_X1  g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G141gat), .ZN(new_n264_));
  INV_X1    g063(.A(G148gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n263_), .A2(KEYINPUT2), .B1(new_n266_), .B2(KEYINPUT3), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n262_), .B(new_n268_), .ZN(new_n269_));
  OAI221_X1 g068(.A(new_n267_), .B1(KEYINPUT3), .B2(new_n266_), .C1(new_n269_), .C2(KEYINPUT2), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT90), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(KEYINPUT1), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n272_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n269_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n266_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G197gat), .B(G204gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT21), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n282_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n286_), .A3(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G228gat), .ZN(new_n289_));
  INV_X1    g088(.A(G233gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n280_), .A2(new_n288_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n280_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n288_), .B(KEYINPUT92), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n261_), .B(new_n293_), .C1(new_n296_), .C2(new_n292_), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n279_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT28), .B1(new_n279_), .B2(KEYINPUT29), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G22gat), .B(G50gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n299_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n300_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n297_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT94), .B(new_n293_), .C1(new_n296_), .C2(new_n292_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT94), .ZN(new_n307_));
  INV_X1    g106(.A(new_n293_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT92), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n288_), .B(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n292_), .B1(new_n310_), .B2(new_n280_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n307_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n261_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT95), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT95), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n306_), .A2(new_n312_), .A3(new_n316_), .A4(new_n313_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n305_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n304_), .A2(new_n301_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(KEYINPUT91), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(KEYINPUT91), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n313_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n320_), .A2(new_n321_), .B1(new_n297_), .B2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT19), .ZN(new_n327_));
  INV_X1    g126(.A(new_n288_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G169gat), .ZN(new_n329_));
  INV_X1    g128(.A(G176gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT84), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n338_), .A2(KEYINPUT85), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(KEYINPUT85), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n334_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n332_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n338_), .A2(new_n336_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  INV_X1    g151(.A(G183gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT25), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G183gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n351_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n344_), .A2(new_n358_), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n325_), .B(new_n327_), .C1(new_n328_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n363_));
  OAI21_X1  g162(.A(G183gat), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT83), .B(G183gat), .C1(new_n362_), .C2(new_n363_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n366_), .A2(new_n355_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n349_), .B1(new_n333_), .B2(new_n346_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n341_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n342_), .B1(new_n338_), .B2(new_n336_), .ZN(new_n371_));
  OAI22_X1  g170(.A1(new_n368_), .A2(new_n370_), .B1(new_n334_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n288_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n372_), .B2(new_n288_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n360_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G8gat), .B(G36gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n288_), .B1(new_n358_), .B2(new_n344_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n384_), .B(KEYINPUT20), .C1(new_n372_), .C2(new_n288_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n327_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n377_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n372_), .A2(new_n288_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT96), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n374_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n392_), .A2(new_n360_), .B1(new_n327_), .B2(new_n385_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(KEYINPUT98), .A3(new_n383_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n377_), .A2(new_n386_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n382_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n389_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT100), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n385_), .A2(new_n327_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n325_), .B1(new_n295_), .B2(new_n359_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n392_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n403_), .B2(new_n327_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT27), .B(new_n387_), .C1(new_n404_), .C2(new_n383_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n399_), .A2(new_n400_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n400_), .B1(new_n399_), .B2(new_n405_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n324_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT101), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412_));
  XOR2_X1   g211(.A(G127gat), .B(G134gat), .Z(new_n413_));
  XOR2_X1   g212(.A(G113gat), .B(G120gat), .Z(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n279_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT99), .ZN(new_n417_));
  INV_X1    g216(.A(new_n415_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n274_), .A2(new_n418_), .A3(new_n278_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n279_), .A2(KEYINPUT99), .A3(new_n415_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n412_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n416_), .A2(KEYINPUT4), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n411_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n410_), .A3(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G85gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT0), .B(G57gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n428_), .B(new_n429_), .Z(new_n430_));
  XNOR2_X1  g229(.A(new_n426_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(G71gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G99gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(G15gat), .B(G43gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT86), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n436_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n372_), .B(KEYINPUT30), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n440_), .A2(KEYINPUT87), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(KEYINPUT87), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n441_), .B2(new_n439_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n415_), .B(KEYINPUT31), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT101), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n324_), .B(new_n450_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n409_), .A2(new_n432_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT88), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n318_), .A2(new_n323_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n383_), .A2(KEYINPUT32), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n393_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n431_), .B(new_n459_), .C1(new_n458_), .C2(new_n404_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n430_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  OR3_X1    g263(.A1(new_n422_), .A2(new_n411_), .A3(new_n423_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n420_), .A2(new_n421_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n430_), .B1(new_n466_), .B2(new_n411_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n397_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n457_), .B1(new_n460_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n399_), .A2(new_n405_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n324_), .A2(new_n431_), .A3(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n456_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n259_), .B1(new_n452_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G230gat), .A2(G233gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT64), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT6), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT6), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  INV_X1    g283(.A(G92gat), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT9), .ZN(new_n486_));
  XOR2_X1   g285(.A(G85gat), .B(G92gat), .Z(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(KEYINPUT9), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT10), .B(G99gat), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n483_), .B(new_n488_), .C1(G106gat), .C2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n478_), .A2(new_n480_), .ZN(new_n492_));
  AND2_X1   g291(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n478_), .B(new_n480_), .C1(new_n494_), .C2(new_n493_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n491_), .B1(new_n502_), .B2(new_n487_), .ZN(new_n503_));
  OR2_X1    g302(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n487_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n483_), .B2(new_n501_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n490_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G71gat), .B(G78gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(KEYINPUT11), .B2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n509_), .A3(KEYINPUT11), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n508_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n490_), .B(new_n515_), .C1(new_n503_), .C2(new_n507_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n517_), .B1(KEYINPUT67), .B2(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(KEYINPUT67), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n476_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n508_), .A2(KEYINPUT68), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n523_), .B(new_n490_), .C1(new_n503_), .C2(new_n507_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n516_), .A2(KEYINPUT12), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n517_), .A2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n518_), .A2(new_n475_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n521_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G120gat), .B(G148gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n521_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(KEYINPUT70), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n540_), .B2(KEYINPUT70), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n539_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n539_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n542_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT72), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n545_), .A2(new_n548_), .B1(new_n549_), .B2(KEYINPUT13), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(KEYINPUT13), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n545_), .A2(new_n548_), .A3(KEYINPUT72), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT78), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n227_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n515_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G127gat), .B(G155gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT16), .ZN(new_n563_));
  XOR2_X1   g362(.A(G183gat), .B(G211gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n561_), .B1(KEYINPUT17), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n565_), .B(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n561_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n508_), .A2(new_n237_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT73), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n522_), .A2(new_n231_), .A3(new_n524_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(new_n581_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT74), .ZN(new_n587_));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(KEYINPUT36), .ZN(new_n591_));
  INV_X1    g390(.A(new_n584_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n576_), .A2(new_n592_), .A3(new_n577_), .A4(new_n582_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n585_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n585_), .B2(new_n593_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n573_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n585_), .A2(new_n593_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n595_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n585_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n572_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n571_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n474_), .A2(new_n557_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(G1gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n431_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n557_), .A2(new_n258_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n571_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n594_), .A2(new_n597_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT102), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n452_), .B2(new_n473_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n432_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n606_), .A2(new_n607_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n608_), .A2(new_n616_), .A3(new_n617_), .ZN(G1324gat));
  NOR2_X1   g417(.A1(new_n406_), .A2(new_n407_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n619_), .A3(new_n610_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G8gat), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT103), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT103), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(KEYINPUT104), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n623_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(G8gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n604_), .A2(new_n629_), .A3(new_n619_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n626_), .A2(KEYINPUT40), .A3(new_n628_), .A4(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n615_), .B2(new_n456_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT41), .Z(new_n637_));
  INV_X1    g436(.A(new_n456_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n604_), .A2(new_n208_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1326gat));
  OAI21_X1  g439(.A(G22gat), .B1(new_n615_), .B2(new_n324_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT42), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n604_), .A2(new_n205_), .A3(new_n457_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1327gat));
  INV_X1    g443(.A(new_n611_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n571_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n474_), .A2(new_n557_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G29gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n431_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n609_), .A2(new_n646_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n452_), .A2(new_n473_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n598_), .A2(new_n602_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n598_), .A2(new_n602_), .ZN(new_n656_));
  AOI211_X1 g455(.A(KEYINPUT43), .B(new_n656_), .C1(new_n452_), .C2(new_n473_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n651_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT44), .B(new_n651_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n431_), .A3(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(KEYINPUT105), .A3(G29gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT105), .B1(new_n662_), .B2(G29gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n650_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n648_), .A2(new_n666_), .A3(new_n619_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT45), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(new_n619_), .A3(new_n661_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(G36gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G36gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI221_X1 g474(.A(new_n668_), .B1(KEYINPUT107), .B2(KEYINPUT46), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  NAND2_X1  g476(.A1(new_n660_), .A2(new_n661_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n449_), .A2(G43gat), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n648_), .A2(new_n638_), .ZN(new_n680_));
  OAI22_X1  g479(.A1(new_n678_), .A2(new_n679_), .B1(G43gat), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g481(.A(G50gat), .B1(new_n678_), .B2(new_n324_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n324_), .A2(G50gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT108), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n648_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1331gat));
  NAND4_X1  g486(.A1(new_n614_), .A2(new_n259_), .A3(new_n556_), .A4(new_n646_), .ZN(new_n688_));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n432_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n258_), .B1(new_n452_), .B2(new_n473_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n556_), .A3(new_n603_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT109), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n432_), .B1(new_n693_), .B2(KEYINPUT110), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(KEYINPUT110), .B2(new_n693_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n690_), .B1(new_n695_), .B2(new_n689_), .ZN(G1332gat));
  INV_X1    g495(.A(new_n619_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G64gat), .B1(new_n688_), .B2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n697_), .A2(G64gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n693_), .B2(new_n701_), .ZN(G1333gat));
  OAI21_X1  g501(.A(G71gat), .B1(new_n688_), .B2(new_n456_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT49), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n638_), .A2(new_n434_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT112), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n693_), .B2(new_n706_), .ZN(G1334gat));
  OAI21_X1  g506(.A(G78gat), .B1(new_n688_), .B2(new_n324_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT50), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n324_), .A2(G78gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n693_), .B2(new_n710_), .ZN(G1335gat));
  AND3_X1   g510(.A1(new_n691_), .A2(new_n556_), .A3(new_n647_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n484_), .A3(new_n431_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n655_), .A2(new_n657_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n557_), .A2(new_n258_), .A3(new_n646_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n431_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n713_), .B1(new_n719_), .B2(new_n484_), .ZN(G1336gat));
  NAND3_X1  g519(.A1(new_n712_), .A2(new_n485_), .A3(new_n619_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n619_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(new_n485_), .ZN(G1337gat));
  OAI21_X1  g523(.A(G99gat), .B1(new_n716_), .B2(new_n456_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n489_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n712_), .A2(new_n449_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g528(.A(new_n715_), .B(new_n457_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT113), .B1(new_n730_), .B2(G106gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT52), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(KEYINPUT52), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G106gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n712_), .A2(new_n736_), .A3(new_n457_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT53), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n733_), .A2(new_n740_), .A3(new_n735_), .A4(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1339gat));
  AND3_X1   g541(.A1(new_n409_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n431_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT59), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n603_), .A2(new_n553_), .A3(new_n259_), .A4(new_n555_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT54), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n527_), .A2(new_n529_), .A3(new_n518_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n476_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n531_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n527_), .A2(new_n529_), .A3(KEYINPUT55), .A4(new_n530_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n538_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n540_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n538_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(KEYINPUT56), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n258_), .A2(new_n756_), .A3(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n246_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT80), .B1(new_n249_), .B2(new_n233_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n240_), .B(new_n255_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n234_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n243_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n255_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n234_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n249_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n254_), .B1(new_n243_), .B2(new_n765_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(KEYINPUT114), .C1(new_n249_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n763_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n760_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n645_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n758_), .A2(KEYINPUT56), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n540_), .A3(new_n756_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n257_), .A2(new_n772_), .A3(new_n770_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT58), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n774_), .A2(new_n784_), .A3(new_n756_), .A4(new_n759_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n654_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n776_), .A2(KEYINPUT57), .A3(new_n645_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n779_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n748_), .B1(new_n646_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n746_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n746_), .A2(KEYINPUT118), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n786_), .B2(new_n654_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT57), .B1(new_n776_), .B2(new_n645_), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n778_), .B(new_n611_), .C1(new_n760_), .C2(new_n775_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n786_), .A2(new_n654_), .A3(new_n797_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n646_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n747_), .B(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n796_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n787_), .A2(KEYINPUT115), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(new_n802_), .A3(new_n779_), .A4(new_n788_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n571_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(KEYINPUT116), .A3(new_n748_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n810_), .A3(new_n744_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(KEYINPUT59), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(KEYINPUT59), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n795_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n258_), .A2(G113gat), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT119), .Z(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n806_), .A2(new_n810_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n258_), .A3(new_n744_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n816_), .A2(new_n818_), .B1(new_n819_), .B2(new_n821_), .ZN(G1340gat));
  OAI21_X1  g621(.A(G120gat), .B1(new_n815_), .B2(new_n557_), .ZN(new_n823_));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n557_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(KEYINPUT60), .B2(new_n824_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n811_), .B2(new_n826_), .ZN(G1341gat));
  OAI21_X1  g626(.A(G127gat), .B1(new_n815_), .B2(new_n571_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n571_), .A2(G127gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n811_), .B2(new_n829_), .ZN(G1342gat));
  NAND2_X1  g629(.A1(new_n654_), .A2(G134gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT120), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n795_), .B(new_n832_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n833_));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n811_), .B2(new_n612_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n838_), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n638_), .A2(new_n324_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n619_), .A2(new_n432_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n806_), .A2(new_n810_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n843_), .A2(new_n844_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n258_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g647(.A(new_n556_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g649(.A(new_n646_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  NOR2_X1   g652(.A1(new_n845_), .A2(new_n846_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G162gat), .B1(new_n854_), .B2(new_n656_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n612_), .A2(G162gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n854_), .B2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(G169gat), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n790_), .A2(new_n324_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n697_), .A2(new_n431_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n638_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n258_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT123), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n858_), .B1(new_n859_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT124), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n866_), .A2(KEYINPUT124), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n859_), .A2(new_n862_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n258_), .A2(new_n329_), .ZN(new_n871_));
  OAI221_X1 g670(.A(new_n869_), .B1(new_n865_), .B2(new_n867_), .C1(new_n870_), .C2(new_n871_), .ZN(G1348gat));
  AND2_X1   g671(.A1(new_n820_), .A2(new_n324_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n861_), .A2(new_n330_), .A3(new_n557_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n859_), .A2(new_n556_), .A3(new_n862_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n873_), .A2(new_n874_), .B1(new_n875_), .B2(new_n330_), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n861_), .A2(new_n571_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G183gat), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n571_), .B(new_n861_), .C1(new_n354_), .C2(new_n357_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n859_), .B2(new_n879_), .ZN(G1350gat));
  OAI21_X1  g679(.A(G190gat), .B1(new_n870_), .B2(new_n656_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n613_), .A2(new_n352_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n870_), .B2(new_n882_), .ZN(G1351gat));
  AND3_X1   g682(.A1(new_n806_), .A2(new_n810_), .A3(new_n841_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n884_), .A2(new_n860_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n258_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n556_), .ZN(new_n888_));
  AND2_X1   g687(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n888_), .B2(new_n889_), .ZN(G1353gat));
  XNOR2_X1  g691(.A(KEYINPUT63), .B(G211gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n885_), .A2(new_n646_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n884_), .A2(new_n860_), .ZN(new_n895_));
  OAI22_X1  g694(.A1(new_n895_), .A2(new_n571_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(new_n899_), .A3(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1354gat));
  OAI21_X1  g700(.A(G218gat), .B1(new_n895_), .B2(new_n656_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n612_), .A2(G218gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n895_), .B2(new_n903_), .ZN(G1355gat));
endmodule


