//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n205_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n204_), .A2(new_n212_), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n214_), .A2(KEYINPUT73), .A3(new_n215_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n213_), .A2(KEYINPUT73), .A3(new_n205_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G229gat), .A3(G233gat), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n204_), .B(KEYINPUT15), .Z(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n212_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n214_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT74), .ZN(new_n226_));
  XOR2_X1   g025(.A(G169gat), .B(G197gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n224_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT6), .Z(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT10), .B(G99gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT64), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(KEYINPUT65), .A3(new_n235_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n232_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT66), .B(G92gat), .Z(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT9), .B1(new_n241_), .B2(G85gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(G85gat), .B2(G92gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G85gat), .B(G92gat), .Z(new_n250_));
  NOR2_X1   g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT7), .Z(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n252_), .B2(new_n232_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT8), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n220_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  OAI221_X1 g057(.A(new_n256_), .B1(KEYINPUT35), .B2(new_n258_), .C1(new_n204_), .C2(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT36), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT103), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT103), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n272_), .A3(new_n269_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n275_), .A2(KEYINPUT1), .A3(G155gat), .A4(G162gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(KEYINPUT84), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n275_), .A2(KEYINPUT1), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT83), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(KEYINPUT82), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n285_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n281_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT85), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n299_), .A3(new_n296_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n284_), .A2(new_n290_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(new_n277_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n294_), .A2(KEYINPUT2), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(KEYINPUT86), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n306_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n305_), .B(new_n307_), .C1(new_n308_), .C2(new_n292_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n298_), .A2(new_n300_), .B1(new_n302_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n301_), .B(new_n277_), .C1(new_n303_), .C2(new_n309_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n291_), .A2(new_n299_), .A3(new_n296_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n299_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT28), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G22gat), .B(G50gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n314_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT91), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT92), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G228gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(G197gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT87), .B1(new_n330_), .B2(G204gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n332_));
  INV_X1    g131(.A(G204gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(G197gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(G204gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT21), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n330_), .B2(G204gat), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n333_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n341_));
  OAI22_X1  g140(.A1(new_n340_), .A2(new_n341_), .B1(new_n330_), .B2(G204gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n337_), .B(new_n338_), .C1(new_n342_), .C2(KEYINPUT21), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT21), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n346_), .B(new_n342_), .C1(new_n345_), .C2(new_n338_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n329_), .B(new_n348_), .C1(new_n311_), .C2(new_n313_), .ZN(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n350_));
  AOI22_X1  g149(.A1(new_n318_), .A2(new_n350_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n329_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n349_), .B(new_n353_), .C1(new_n329_), .C2(new_n351_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n323_), .A2(KEYINPUT91), .A3(new_n324_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n325_), .A2(new_n326_), .A3(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n328_), .A2(new_n357_), .A3(new_n358_), .A4(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n363_));
  AOI211_X1 g162(.A(KEYINPUT91), .B(KEYINPUT92), .C1(new_n323_), .C2(new_n324_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT101), .ZN(new_n368_));
  XOR2_X1   g167(.A(G8gat), .B(G36gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT100), .Z(new_n373_));
  NOR2_X1   g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G169gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n382_));
  INV_X1    g181(.A(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(G176gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT24), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n376_), .B(KEYINPUT23), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT25), .B(G183gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n388_), .B1(G169gat), .B2(G176gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .A4(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n343_), .A2(new_n347_), .A3(new_n381_), .A4(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT98), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n389_), .A2(KEYINPUT76), .A3(new_n390_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT24), .B1(new_n385_), .B2(new_n386_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n376_), .B(new_n375_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n401_), .A2(new_n405_), .A3(new_n393_), .A4(new_n395_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n378_), .A2(KEYINPUT77), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n374_), .A2(KEYINPUT77), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n390_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(new_n380_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n406_), .A2(new_n410_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT98), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n397_), .A2(new_n413_), .A3(new_n398_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n400_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT19), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n396_), .A2(new_n381_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n348_), .B2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n406_), .A2(new_n410_), .A3(new_n343_), .A4(new_n347_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n417_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n373_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n397_), .A2(KEYINPUT20), .A3(new_n423_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n428_), .A2(new_n411_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n429_), .A3(new_n372_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT27), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n368_), .B1(new_n425_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n428_), .A2(new_n411_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n426_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n433_), .B1(new_n435_), .B2(new_n372_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n424_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n436_), .B(KEYINPUT101), .C1(new_n438_), .C2(new_n373_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n372_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n426_), .B2(new_n434_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n430_), .A2(new_n441_), .A3(KEYINPUT93), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n427_), .A2(new_n429_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT93), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n440_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n433_), .A3(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n432_), .A2(new_n439_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n367_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT96), .ZN(new_n450_));
  XOR2_X1   g249(.A(G127gat), .B(G134gat), .Z(new_n451_));
  XOR2_X1   g250(.A(G113gat), .B(G120gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n318_), .A2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n453_), .B(new_n315_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT94), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT94), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n318_), .A2(new_n458_), .A3(new_n454_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n450_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  AOI211_X1 g262(.A(KEYINPUT96), .B(new_n463_), .C1(new_n457_), .C2(new_n459_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT4), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n298_), .A2(new_n300_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n453_), .B1(new_n467_), .B2(new_n315_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n465_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n463_), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n462_), .A2(new_n464_), .B1(new_n466_), .B2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G1gat), .B(G29gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n462_), .A2(new_n464_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT99), .ZN(new_n479_));
  INV_X1    g278(.A(new_n476_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n466_), .B2(new_n470_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n456_), .A2(KEYINPUT94), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(new_n468_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n459_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n461_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT96), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n460_), .A2(new_n450_), .A3(new_n461_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n460_), .A2(KEYINPUT4), .ZN(new_n490_));
  INV_X1    g289(.A(new_n470_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n476_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT99), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n477_), .B1(new_n482_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n406_), .A2(new_n410_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G227gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G15gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n495_), .B(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G71gat), .B(G99gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT79), .B(G43gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n498_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n453_), .B(KEYINPUT31), .Z(new_n507_));
  OR2_X1    g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n505_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n509_), .A3(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n494_), .A2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n449_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n511_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n438_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n372_), .A2(KEYINPUT32), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n443_), .B2(new_n516_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n479_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n489_), .A2(KEYINPUT99), .A3(new_n492_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n521_), .B2(new_n477_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT33), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n489_), .A2(KEYINPUT33), .A3(new_n492_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n490_), .A2(new_n461_), .A3(new_n469_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n480_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n526_), .A2(new_n527_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n366_), .B1(new_n522_), .B2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n447_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n519_), .A2(new_n520_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n514_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n513_), .B1(new_n535_), .B2(KEYINPUT102), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT102), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n529_), .B1(new_n533_), .B2(new_n518_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n538_), .A2(new_n366_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(new_n514_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n274_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(G230gat), .ZN(new_n542_));
  INV_X1    g341(.A(G233gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n253_), .B(KEYINPUT8), .Z(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n240_), .B2(new_n248_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT68), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G78gat), .Z(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(KEYINPUT11), .B2(new_n548_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n550_), .B(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n546_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n249_), .A2(new_n553_), .A3(new_n254_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT69), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n546_), .A2(new_n553_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n544_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n544_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n546_), .A2(KEYINPUT12), .A3(new_n553_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(new_n553_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n255_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n560_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT5), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n559_), .A2(new_n565_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT13), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(KEYINPUT70), .B2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n212_), .B(KEYINPUT71), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n563_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT72), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n583_), .A2(new_n592_), .A3(new_n587_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT72), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND4_X1   g395(.A1(new_n230_), .A2(new_n541_), .A3(new_n579_), .A4(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n597_), .A2(new_n494_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n207_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n229_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n270_), .A2(KEYINPUT37), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n267_), .A2(new_n603_), .A3(new_n269_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n595_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n601_), .A2(new_n579_), .A3(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n207_), .A3(new_n494_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n599_), .B1(new_n600_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n600_), .B2(new_n609_), .ZN(G1324gat));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n208_), .A3(new_n448_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n597_), .A2(new_n448_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n614_), .B2(G8gat), .ZN(new_n615_));
  AOI211_X1 g414(.A(KEYINPUT39), .B(new_n208_), .C1(new_n597_), .C2(new_n448_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT40), .B(new_n612_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1325gat));
  INV_X1    g420(.A(G15gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n597_), .B2(new_n514_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT41), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n608_), .A2(new_n622_), .A3(new_n514_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1326gat));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n608_), .A2(new_n627_), .A3(new_n367_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n597_), .A2(new_n367_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G22gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT105), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n632_), .A3(G22gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n634_));
  AND3_X1   g433(.A1(new_n631_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n628_), .B1(new_n635_), .B2(new_n636_), .ZN(G1327gat));
  AND4_X1   g436(.A1(new_n601_), .A2(new_n579_), .A3(new_n595_), .A4(new_n274_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G29gat), .B1(new_n638_), .B2(new_n494_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n579_), .A2(new_n230_), .A3(new_n595_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI211_X1 g440(.A(KEYINPUT43), .B(new_n605_), .C1(new_n536_), .C2(new_n540_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n513_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n518_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n494_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n367_), .B1(new_n647_), .B2(new_n529_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n494_), .A2(new_n366_), .A3(new_n448_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT102), .B(new_n511_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n540_), .A2(new_n645_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n644_), .B1(new_n651_), .B2(new_n606_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT44), .B(new_n641_), .C1(new_n642_), .C2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT107), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n655_), .A3(new_n606_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n605_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n644_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(KEYINPUT44), .A4(new_n641_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n654_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n641_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n494_), .A2(G29gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n639_), .B1(new_n665_), .B2(new_n666_), .ZN(G1328gat));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(KEYINPUT46), .ZN(new_n669_));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n662_), .A2(new_n447_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n661_), .B2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n447_), .A2(G36gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n638_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n669_), .B1(new_n672_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n669_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n651_), .A2(new_n606_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n643_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n640_), .B1(new_n681_), .B2(new_n656_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n448_), .B1(new_n682_), .B2(KEYINPUT44), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n654_), .B2(new_n660_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n678_), .B(new_n679_), .C1(new_n684_), .C2(new_n670_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n677_), .A2(new_n685_), .ZN(G1329gat));
  NAND2_X1  g485(.A1(new_n514_), .A2(G43gat), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n687_), .B(new_n662_), .C1(new_n654_), .C2(new_n660_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n638_), .A2(new_n514_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(G43gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT47), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  INV_X1    g491(.A(new_n690_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n692_), .B(new_n693_), .C1(new_n664_), .C2(new_n687_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1330gat));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n638_), .A2(new_n696_), .A3(new_n367_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n658_), .A2(new_n641_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n366_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n661_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n698_), .B1(new_n702_), .B2(G50gat), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT109), .B(new_n696_), .C1(new_n661_), .C2(new_n701_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n697_), .B1(new_n703_), .B2(new_n704_), .ZN(G1331gat));
  AOI21_X1  g504(.A(new_n230_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n579_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n607_), .ZN(new_n708_));
  INV_X1    g507(.A(G57gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n494_), .ZN(new_n710_));
  AND4_X1   g509(.A1(new_n229_), .A2(new_n541_), .A3(new_n707_), .A4(new_n596_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n494_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n712_), .B2(new_n709_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n711_), .B2(new_n448_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n708_), .A2(new_n714_), .A3(new_n448_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n711_), .B2(new_n514_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT49), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n708_), .A2(new_n720_), .A3(new_n514_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1334gat));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n711_), .B2(new_n367_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT50), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n708_), .A2(new_n725_), .A3(new_n367_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1335gat));
  INV_X1    g528(.A(new_n274_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n730_), .A2(new_n579_), .A3(new_n596_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n706_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(G85gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n494_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n579_), .A2(new_n230_), .A3(new_n596_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT111), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n658_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n494_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n739_), .B2(new_n733_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n732_), .B2(new_n448_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n448_), .A2(new_n241_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n737_), .B2(new_n742_), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n732_), .A2(new_n514_), .A3(new_n234_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT112), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n737_), .A2(new_n514_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G99gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n745_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n732_), .A2(new_n235_), .A3(new_n367_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n658_), .A2(new_n736_), .A3(new_n367_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(G106gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G106gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n752_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  NAND2_X1  g560(.A1(new_n230_), .A2(new_n571_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n560_), .B(KEYINPUT55), .C1(new_n561_), .C2(new_n564_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT117), .ZN(new_n764_));
  INV_X1    g563(.A(new_n544_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n555_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT12), .B1(new_n546_), .B2(new_n553_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n255_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(KEYINPUT55), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n556_), .B(new_n554_), .C1(new_n561_), .C2(new_n564_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n772_), .A2(KEYINPUT116), .A3(new_n544_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT116), .B1(new_n772_), .B2(new_n544_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n764_), .B(new_n771_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n769_), .B2(KEYINPUT55), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n565_), .A2(KEYINPUT115), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n569_), .B1(new_n775_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT118), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n764_), .A2(new_n771_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(new_n780_), .C1(new_n774_), .C2(new_n773_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(new_n569_), .A3(new_n784_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n762_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n219_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n218_), .A2(new_n222_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n222_), .B1(new_n205_), .B2(new_n213_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n228_), .B1(new_n221_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(new_n792_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n791_), .A2(new_n796_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n574_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n730_), .B1(new_n790_), .B2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n762_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n789_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n784_), .B1(new_n788_), .B2(new_n569_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n800_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n802_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n730_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n803_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n788_), .A2(new_n783_), .A3(new_n569_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n799_), .A2(new_n797_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n571_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT121), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n818_), .A3(new_n571_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n814_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n783_), .B1(new_n788_), .B2(new_n569_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n813_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n606_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(KEYINPUT58), .A3(new_n814_), .A4(new_n820_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n827_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n595_), .B1(new_n812_), .B2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n605_), .A2(new_n579_), .A3(new_n229_), .A4(new_n596_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n833_));
  AND2_X1   g632(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n833_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n449_), .A2(new_n514_), .A3(new_n494_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT123), .Z(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n230_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n839_), .A2(KEYINPUT59), .A3(new_n841_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n229_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n849_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n579_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n843_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n579_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n843_), .B2(new_n596_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n847_), .A2(new_n848_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n595_), .A2(KEYINPUT124), .ZN(new_n858_));
  MUX2_X1   g657(.A(KEYINPUT124), .B(new_n858_), .S(G127gat), .Z(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n857_), .B2(new_n859_), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n843_), .A2(new_n861_), .A3(new_n274_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n605_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n514_), .A2(new_n533_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n839_), .A2(new_n532_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n229_), .ZN(new_n867_));
  INV_X1    g666(.A(G141gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n579_), .ZN(new_n870_));
  INV_X1    g669(.A(G148gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n866_), .A2(new_n595_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n866_), .B2(new_n605_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n730_), .A2(G162gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n866_), .B2(new_n877_), .ZN(G1347gat));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(KEYINPUT125), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n367_), .A2(new_n494_), .A3(new_n511_), .A4(new_n447_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n839_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(G169gat), .B(new_n880_), .C1(new_n882_), .C2(new_n229_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n882_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT22), .B(G169gat), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n230_), .A2(new_n885_), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(KEYINPUT126), .Z(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n383_), .B1(new_n884_), .B2(new_n230_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n890_));
  OAI211_X1 g689(.A(new_n883_), .B(new_n888_), .C1(new_n889_), .C2(new_n890_), .ZN(G1348gat));
  NOR2_X1   g690(.A1(new_n882_), .A2(new_n579_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n384_), .ZN(G1349gat));
  AOI21_X1  g692(.A(G183gat), .B1(new_n884_), .B2(new_n596_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n882_), .A2(new_n391_), .A3(new_n595_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n882_), .B2(new_n605_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n274_), .A2(new_n392_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n882_), .B2(new_n898_), .ZN(G1351gat));
  INV_X1    g698(.A(KEYINPUT127), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n825_), .A2(new_n814_), .A3(new_n820_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n605_), .B1(new_n901_), .B2(new_n813_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n826_), .A2(new_n827_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n826_), .A2(new_n827_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n811_), .A3(new_n803_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n837_), .B1(new_n906_), .B2(new_n595_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n514_), .A2(new_n494_), .A3(new_n366_), .A4(new_n447_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n900_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n810_), .B1(new_n809_), .B2(new_n730_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n274_), .B(new_n802_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n596_), .B1(new_n913_), .B2(new_n905_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT127), .B(new_n908_), .C1(new_n914_), .C2(new_n837_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n910_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916_), .B2(new_n230_), .ZN(new_n917_));
  AOI211_X1 g716(.A(new_n330_), .B(new_n229_), .C1(new_n910_), .C2(new_n915_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1352gat));
  AOI21_X1  g718(.A(KEYINPUT127), .B1(new_n839_), .B2(new_n908_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n907_), .A2(new_n900_), .A3(new_n909_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n707_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(G204gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n916_), .A2(new_n333_), .A3(new_n707_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1353gat));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n595_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n916_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n928_), .ZN(new_n930_));
  AOI211_X1 g729(.A(new_n926_), .B(new_n930_), .C1(new_n910_), .C2(new_n915_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1354gat));
  INV_X1    g731(.A(G218gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n916_), .A2(new_n933_), .A3(new_n274_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n605_), .B1(new_n910_), .B2(new_n915_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n933_), .B2(new_n935_), .ZN(G1355gat));
endmodule


