//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G64gat), .B(G92gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT99), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT100), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G8gat), .B(G36gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT106), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G226gat), .A2(G233gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT19), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT20), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT91), .ZN(new_n215_));
  INV_X1    g014(.A(G211gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(G218gat), .ZN(new_n217_));
  INV_X1    g016(.A(G218gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(G211gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n215_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(G211gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(G218gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT91), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(G204gat), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(KEYINPUT21), .A3(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n232_));
  INV_X1    g031(.A(G197gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(G204gat), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT90), .ZN(new_n237_));
  INV_X1    g036(.A(G204gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(G197gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT21), .B1(new_n236_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n238_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n228_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n245_), .A3(new_n224_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT92), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n227_), .A2(new_n229_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n249_), .A2(new_n243_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(KEYINPUT92), .A3(new_n242_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n231_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT23), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT23), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(G183gat), .A3(G190gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT81), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT81), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n253_), .B2(KEYINPUT23), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n257_), .A2(new_n259_), .B1(G183gat), .B2(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(G169gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT22), .B1(new_n261_), .B2(KEYINPUT79), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(G169gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(KEYINPUT80), .A2(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(KEYINPUT80), .A2(G176gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n262_), .A2(new_n265_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G176gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n261_), .A2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n272_), .A2(KEYINPUT24), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(KEYINPUT24), .A3(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT25), .B(G183gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G190gat), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n277_), .A2(new_n278_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n260_), .A2(new_n270_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n214_), .B1(new_n252_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT97), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n254_), .A2(new_n256_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(G183gat), .B2(G190gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT22), .B(G169gat), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n266_), .A2(new_n267_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(G169gat), .B2(G176gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n257_), .A2(new_n259_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(new_n275_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n278_), .A2(KEYINPUT96), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n278_), .A2(KEYINPUT96), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n277_), .A3(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n284_), .A2(new_n288_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n252_), .A2(new_n282_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n231_), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT92), .B1(new_n250_), .B2(new_n242_), .ZN(new_n297_));
  AND4_X1   g096(.A1(KEYINPUT92), .A2(new_n242_), .A3(new_n245_), .A4(new_n224_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n288_), .A2(new_n284_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n290_), .A2(new_n293_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT97), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n213_), .B(new_n281_), .C1(new_n295_), .C2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n270_), .A2(new_n260_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n276_), .A2(new_n279_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n299_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n252_), .A2(new_n294_), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT105), .B(KEYINPUT20), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n212_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n210_), .B1(new_n304_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT20), .B1(new_n299_), .B2(new_n307_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n282_), .B1(new_n252_), .B2(new_n294_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n299_), .A2(KEYINPUT97), .A3(new_n302_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT106), .B1(new_n318_), .B2(new_n213_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n209_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT108), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT108), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n209_), .C1(new_n314_), .C2(new_n319_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n209_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n212_), .A2(new_n214_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n308_), .A2(new_n309_), .A3(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n324_), .B(new_n326_), .C1(new_n318_), .C2(new_n213_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n321_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT27), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n316_), .A2(new_n317_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n213_), .B1(new_n330_), .B2(new_n281_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n326_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n209_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(KEYINPUT101), .A3(new_n327_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n281_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(new_n212_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT101), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n324_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT27), .B1(new_n334_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT86), .ZN(new_n347_));
  OAI221_X1 g146(.A(new_n347_), .B1(KEYINPUT85), .B2(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT87), .B(KEYINPUT2), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT2), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n353_), .A2(new_n350_), .B1(KEYINPUT86), .B2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(KEYINPUT86), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n351_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT84), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT83), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT84), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n361_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n361_), .B(KEYINPUT1), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n365_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n366_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n350_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(new_n356_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  OAI22_X1  g177(.A1(new_n360_), .A2(new_n369_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT88), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(KEYINPUT87), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n352_), .A2(KEYINPUT2), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n376_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(new_n358_), .A3(new_n355_), .A4(new_n348_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n373_), .A2(new_n374_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n361_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n361_), .B(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n377_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n392_), .A3(KEYINPUT88), .ZN(new_n393_));
  XOR2_X1   g192(.A(G127gat), .B(G134gat), .Z(new_n394_));
  XOR2_X1   g193(.A(G113gat), .B(G120gat), .Z(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  NAND3_X1  g195(.A1(new_n381_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n379_), .A2(new_n396_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n346_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n388_), .A2(new_n392_), .A3(KEYINPUT88), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT88), .B1(new_n388_), .B2(new_n392_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT4), .B1(new_n403_), .B2(new_n396_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n400_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n398_), .B1(new_n403_), .B2(new_n396_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n405_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n345_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT107), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n397_), .A2(new_n346_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n408_), .B(new_n412_), .C1(new_n407_), .C2(new_n346_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n407_), .A2(new_n408_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n345_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n410_), .A2(new_n411_), .A3(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT107), .B(new_n345_), .C1(new_n406_), .C2(new_n409_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(G15gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT30), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT31), .ZN(new_n425_));
  INV_X1    g224(.A(new_n396_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G43gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n307_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n280_), .A2(new_n428_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n426_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n431_), .A3(new_n426_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n425_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n434_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n425_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n432_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT82), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n435_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(G228gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n299_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n248_), .A2(new_n251_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n445_), .B1(new_n450_), .B2(new_n296_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n381_), .A2(KEYINPUT29), .A3(new_n393_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n445_), .A2(new_n449_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G78gat), .B(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT94), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n451_), .A2(new_n452_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n445_), .B1(new_n252_), .B2(new_n447_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n455_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(KEYINPUT95), .A3(new_n455_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n456_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT95), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G22gat), .B(G50gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n446_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT28), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT28), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n470_), .B(new_n446_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n471_), .A3(new_n467_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n463_), .A2(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n469_), .A2(new_n471_), .A3(new_n467_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(new_n472_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n464_), .A2(KEYINPUT93), .ZN(new_n479_));
  INV_X1    g278(.A(new_n459_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n457_), .A2(new_n458_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT93), .A3(new_n454_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n478_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n444_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n460_), .B1(new_n482_), .B2(new_n454_), .ZN(new_n486_));
  AND4_X1   g285(.A1(KEYINPUT95), .A2(new_n457_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n478_), .A3(new_n466_), .A4(new_n461_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n459_), .B1(KEYINPUT93), .B2(new_n464_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n483_), .ZN(new_n491_));
  OAI22_X1  g290(.A1(new_n490_), .A2(new_n491_), .B1(new_n477_), .B2(new_n472_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n435_), .A2(new_n439_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n420_), .B1(new_n485_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n415_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT33), .B1(new_n496_), .B2(KEYINPUT102), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT102), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n410_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n345_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n412_), .B1(new_n407_), .B2(new_n346_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT103), .B1(new_n502_), .B2(new_n405_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT103), .B(new_n405_), .C1(new_n400_), .C2(new_n404_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n501_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(new_n500_), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n334_), .A2(new_n338_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n336_), .B2(KEYINPUT104), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n314_), .A2(new_n319_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT104), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n336_), .A2(new_n512_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n510_), .A2(new_n511_), .B1(new_n513_), .B2(new_n509_), .ZN(new_n514_));
  OAI22_X1  g313(.A1(new_n507_), .A2(new_n508_), .B1(new_n514_), .B2(new_n419_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n489_), .A2(new_n492_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n444_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n341_), .A2(new_n495_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G190gat), .B(G218gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G134gat), .B(G162gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(KEYINPUT36), .Z(new_n523_));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G232gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT34), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528_));
  XOR2_X1   g327(.A(G29gat), .B(G36gat), .Z(new_n529_));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G29gat), .B(G36gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT72), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n528_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n533_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(KEYINPUT15), .A3(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G99gat), .ZN(new_n544_));
  INV_X1    g343(.A(G106gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT6), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(G99gat), .A3(G106gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT64), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT7), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n550_), .A2(new_n553_), .A3(new_n544_), .A4(new_n545_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G85gat), .B(G92gat), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(KEYINPUT65), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT66), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(KEYINPUT66), .A3(new_n556_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n559_), .A2(KEYINPUT8), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT8), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT10), .B(G99gat), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n545_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n556_), .A2(KEYINPUT9), .ZN(new_n566_));
  INV_X1    g365(.A(G85gat), .ZN(new_n567_));
  INV_X1    g366(.A(G92gat), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n567_), .A2(new_n568_), .A3(KEYINPUT9), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n565_), .A2(new_n566_), .A3(new_n549_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n543_), .B1(new_n561_), .B2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n563_), .A2(new_n570_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n540_), .A2(new_n541_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n559_), .A2(KEYINPUT8), .A3(new_n560_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n524_), .B(new_n527_), .C1(new_n572_), .C2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n527_), .A2(new_n524_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n527_), .A2(new_n524_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n572_), .A2(new_n579_), .A3(new_n580_), .A4(new_n576_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n523_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n537_), .A2(new_n542_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n578_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n522_), .A2(KEYINPUT36), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n581_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n519_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT68), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT11), .ZN(new_n594_));
  XOR2_X1   g393(.A(G71gat), .B(G78gat), .Z(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n593_), .A2(KEYINPUT11), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n595_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n601_));
  OAI21_X1  g400(.A(new_n592_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n573_), .A2(new_n575_), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n599_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n606_), .B1(new_n561_), .B2(new_n571_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n601_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(KEYINPUT68), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n600_), .A2(KEYINPUT12), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n602_), .A2(new_n605_), .A3(new_n609_), .A4(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n603_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(G230gat), .A3(G233gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(G120gat), .B(G148gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT70), .ZN(new_n615_));
  XOR2_X1   g414(.A(G176gat), .B(G204gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n611_), .A2(new_n613_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT71), .ZN(new_n622_));
  OAI22_X1  g421(.A1(new_n620_), .A2(new_n621_), .B1(new_n622_), .B2(KEYINPUT13), .ZN(new_n623_));
  INV_X1    g422(.A(new_n621_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n611_), .A2(new_n613_), .A3(new_n619_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(G8gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT74), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT74), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n632_), .B(KEYINPUT14), .C1(new_n202_), .C2(new_n629_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G15gat), .B(G22gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G1gat), .B(G8gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n635_), .B(new_n636_), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(new_n574_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G229gat), .A2(G233gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n637_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n543_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n637_), .A2(new_n574_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n639_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT78), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n646_), .B(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n628_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(G231gat), .A2(G233gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n599_), .B(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT75), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(new_n637_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT77), .ZN(new_n660_));
  XNOR2_X1  g459(.A(G127gat), .B(G155gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(G183gat), .B(G211gat), .Z(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT17), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n657_), .B(new_n642_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n664_), .B(KEYINPUT17), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n654_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n591_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n202_), .B1(new_n673_), .B2(new_n420_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT110), .Z(new_n675_));
  NOR2_X1   g474(.A1(new_n519_), .A2(new_n652_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n583_), .A2(new_n589_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n583_), .A2(KEYINPUT73), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(KEYINPUT37), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT37), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n583_), .B(new_n589_), .C1(KEYINPUT73), .C2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n671_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n628_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n202_), .A2(new_n676_), .A3(new_n420_), .A4(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(KEYINPUT38), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT111), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(KEYINPUT38), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT109), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n675_), .A2(new_n688_), .A3(new_n690_), .ZN(G1324gat));
  AND2_X1   g490(.A1(new_n676_), .A2(new_n685_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n341_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n629_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n591_), .A2(new_n693_), .A3(new_n672_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT39), .ZN(new_n697_));
  AND4_X1   g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .A4(G8gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n629_), .B1(KEYINPUT112), .B2(KEYINPUT39), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n696_), .A2(new_n699_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n694_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1325gat));
  NAND2_X1  g502(.A1(new_n673_), .A2(new_n517_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G15gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT113), .B(KEYINPUT41), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n692_), .A2(new_n422_), .A3(new_n517_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(G1326gat));
  INV_X1    g509(.A(G22gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n673_), .B2(new_n516_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT42), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n692_), .A2(new_n711_), .A3(new_n516_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1327gat));
  INV_X1    g514(.A(KEYINPUT114), .ZN(new_n716_));
  INV_X1    g515(.A(new_n523_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n587_), .B2(new_n581_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT73), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT37), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n590_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n681_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n716_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n679_), .A2(KEYINPUT114), .A3(new_n681_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n485_), .A2(new_n494_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT27), .ZN(new_n727_));
  INV_X1    g526(.A(new_n327_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n320_), .B2(KEYINPUT108), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n729_), .B2(new_n323_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n419_), .B(new_n726_), .C1(new_n730_), .C2(new_n339_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n515_), .A2(new_n518_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n725_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n679_), .A2(new_n681_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n734_), .ZN(new_n737_));
  OAI22_X1  g536(.A1(new_n733_), .A2(new_n734_), .B1(new_n519_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n671_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n654_), .A2(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n738_), .A2(KEYINPUT44), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT44), .B1(new_n738_), .B2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n420_), .A2(G29gat), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n671_), .A2(new_n590_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n684_), .A2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n676_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G29gat), .B1(new_n747_), .B2(new_n420_), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n744_), .A2(KEYINPUT115), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT115), .B1(new_n744_), .B2(new_n748_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1328gat));
  INV_X1    g550(.A(G36gat), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n676_), .A2(new_n752_), .A3(new_n693_), .A4(new_n746_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT45), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n741_), .A2(new_n742_), .A3(new_n341_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n752_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT46), .B(new_n754_), .C1(new_n755_), .C2(new_n752_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1329gat));
  NAND2_X1  g559(.A1(new_n493_), .A2(G43gat), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n741_), .A2(new_n742_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G43gat), .B1(new_n747_), .B2(new_n517_), .ZN(new_n763_));
  OR3_X1    g562(.A1(new_n762_), .A2(KEYINPUT47), .A3(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT47), .B1(new_n762_), .B2(new_n763_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1330gat));
  AOI21_X1  g565(.A(G50gat), .B1(new_n747_), .B2(new_n516_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n741_), .A2(new_n742_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n516_), .A2(G50gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(G1331gat));
  NOR4_X1   g569(.A1(new_n519_), .A2(new_n653_), .A3(new_n628_), .A4(new_n683_), .ZN(new_n771_));
  INV_X1    g570(.A(G57gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n420_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n684_), .A2(new_n652_), .ZN(new_n774_));
  NOR4_X1   g573(.A1(new_n519_), .A2(new_n590_), .A3(new_n671_), .A4(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(new_n420_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n773_), .B1(new_n776_), .B2(new_n772_), .ZN(G1332gat));
  INV_X1    g576(.A(G64gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n775_), .B2(new_n693_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT48), .Z(new_n780_));
  NAND3_X1  g579(.A1(new_n771_), .A2(new_n778_), .A3(new_n693_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1333gat));
  INV_X1    g581(.A(G71gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n775_), .B2(new_n517_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT49), .Z(new_n785_));
  NAND3_X1  g584(.A1(new_n771_), .A2(new_n783_), .A3(new_n517_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1334gat));
  INV_X1    g586(.A(G78gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n771_), .A2(new_n788_), .A3(new_n516_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n775_), .B2(new_n516_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(new_n791_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(G1335gat));
  NOR2_X1   g593(.A1(new_n774_), .A2(new_n739_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n738_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n419_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n519_), .A2(new_n653_), .A3(new_n628_), .A4(new_n745_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n567_), .A3(new_n420_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1336gat));
  OAI21_X1  g599(.A(G92gat), .B1(new_n796_), .B2(new_n341_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n568_), .A3(new_n693_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n796_), .B2(new_n444_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n493_), .A2(new_n564_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n798_), .A2(new_n805_), .B1(new_n806_), .B2(KEYINPUT51), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(KEYINPUT51), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n808_), .B(new_n809_), .Z(G1338gat));
  NAND3_X1  g609(.A1(new_n798_), .A2(new_n545_), .A3(new_n516_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n738_), .A2(new_n516_), .A3(new_n795_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(G106gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n812_), .B2(G106gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT53), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n811_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1339gat));
  INV_X1    g619(.A(new_n494_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n341_), .A2(new_n420_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n638_), .A2(new_n639_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n643_), .A2(new_n644_), .A3(new_n640_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n650_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n823_), .A2(new_n824_), .A3(KEYINPUT120), .A4(new_n650_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n646_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n827_), .A2(new_n828_), .B1(new_n829_), .B2(new_n649_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n625_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n602_), .A2(new_n609_), .A3(new_n603_), .A4(new_n610_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(G230gat), .A3(G233gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n573_), .A2(new_n575_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n601_), .B1(new_n834_), .B2(new_n606_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n835_), .A2(KEYINPUT68), .B1(KEYINPUT12), .B2(new_n600_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT55), .A3(new_n602_), .A4(new_n605_), .ZN(new_n837_));
  XOR2_X1   g636(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n838_));
  NAND2_X1  g637(.A1(new_n611_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n833_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n619_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n841_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n831_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n736_), .B1(new_n846_), .B2(KEYINPUT58), .ZN(new_n847_));
  INV_X1    g646(.A(new_n831_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n841_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n841_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT58), .B(new_n848_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n620_), .A2(new_n652_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n626_), .A2(new_n830_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n590_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n847_), .A2(new_n852_), .B1(new_n856_), .B2(KEYINPUT57), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(KEYINPUT57), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n671_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n628_), .A2(new_n735_), .A3(new_n739_), .A4(new_n652_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT118), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n682_), .A2(new_n863_), .A3(new_n652_), .A4(new_n628_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(KEYINPUT54), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT54), .B1(new_n862_), .B2(new_n864_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n822_), .B1(new_n860_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G113gat), .B1(new_n869_), .B2(new_n653_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  INV_X1    g670(.A(new_n822_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873_));
  INV_X1    g672(.A(new_n853_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n855_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n677_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n735_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n873_), .A2(new_n877_), .B1(new_n880_), .B2(new_n851_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n739_), .B1(new_n881_), .B2(new_n858_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n862_), .A2(new_n864_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n865_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n871_), .B(new_n872_), .C1(new_n882_), .C2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n881_), .A2(new_n858_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n886_), .B1(new_n671_), .B2(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n892_), .C2(new_n822_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n888_), .B1(new_n890_), .B2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n653_), .A2(KEYINPUT122), .A3(G113gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(KEYINPUT122), .B2(G113gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n870_), .B1(new_n894_), .B2(new_n896_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n628_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n869_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n887_), .A2(new_n684_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n890_), .B2(new_n893_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n902_), .B2(new_n898_), .ZN(G1341gat));
  AOI21_X1  g702(.A(G127gat), .B1(new_n869_), .B2(new_n739_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n739_), .A2(G127gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT123), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n894_), .B2(new_n906_), .ZN(G1342gat));
  AOI21_X1  g706(.A(G134gat), .B1(new_n869_), .B2(new_n590_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT124), .B(G134gat), .Z(new_n909_));
  NOR2_X1   g708(.A1(new_n735_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n894_), .B2(new_n910_), .ZN(G1343gat));
  NAND2_X1  g710(.A1(new_n860_), .A2(new_n868_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n693_), .A2(new_n419_), .A3(new_n485_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n653_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(G141gat), .ZN(new_n916_));
  INV_X1    g715(.A(G141gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n917_), .A3(new_n653_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n684_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G148gat), .ZN(new_n921_));
  INV_X1    g720(.A(G148gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n914_), .A2(new_n922_), .A3(new_n684_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1345gat));
  OAI211_X1 g723(.A(new_n739_), .B(new_n913_), .C1(new_n882_), .C2(new_n886_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT125), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n912_), .A2(new_n927_), .A3(new_n739_), .A4(new_n913_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT61), .B(G155gat), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n926_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1346gat));
  AOI21_X1  g731(.A(G162gat), .B1(new_n914_), .B2(new_n590_), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n723_), .A2(G162gat), .A3(new_n724_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n914_), .B2(new_n934_), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n341_), .A2(new_n420_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n516_), .A2(new_n444_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n912_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G169gat), .B1(new_n938_), .B2(new_n652_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  OR3_X1    g740(.A1(new_n938_), .A2(new_n285_), .A3(new_n652_), .ZN(new_n942_));
  OAI211_X1 g741(.A(KEYINPUT62), .B(G169gat), .C1(new_n938_), .C2(new_n652_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(G1348gat));
  NOR2_X1   g743(.A1(new_n938_), .A2(new_n628_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n286_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n938_), .A2(new_n271_), .A3(new_n628_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1349gat));
  NOR2_X1   g747(.A1(new_n938_), .A2(new_n671_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(G183gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n938_), .A2(new_n277_), .A3(new_n671_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n938_), .B2(new_n735_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n590_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n938_), .B2(new_n954_), .ZN(G1351gat));
  INV_X1    g754(.A(new_n485_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n912_), .A2(new_n956_), .A3(new_n936_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n233_), .A2(KEYINPUT126), .ZN(new_n958_));
  OR3_X1    g757(.A1(new_n957_), .A2(new_n652_), .A3(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n233_), .A2(KEYINPUT126), .ZN(new_n960_));
  OAI22_X1  g759(.A1(new_n957_), .A2(new_n652_), .B1(new_n960_), .B2(new_n958_), .ZN(new_n961_));
  AND2_X1   g760(.A1(new_n959_), .A2(new_n961_), .ZN(G1352gat));
  NOR2_X1   g761(.A1(new_n957_), .A2(new_n628_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(new_n238_), .ZN(G1353gat));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n739_), .B1(new_n965_), .B2(new_n216_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n957_), .A2(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n216_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(KEYINPUT127), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n967_), .B(new_n969_), .ZN(G1354gat));
  OAI21_X1  g769(.A(G218gat), .B1(new_n957_), .B2(new_n735_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n590_), .A2(new_n218_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n957_), .B2(new_n972_), .ZN(G1355gat));
endmodule


