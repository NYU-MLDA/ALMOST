//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_;
  AND2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT64), .B1(new_n202_), .B2(KEYINPUT9), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(new_n202_), .B2(KEYINPUT9), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT65), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n213_), .A3(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT10), .B(G99gat), .Z(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n212_), .A2(new_n214_), .A3(new_n219_), .A4(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n202_), .B2(new_n209_), .ZN(new_n229_));
  INV_X1    g028(.A(G85gat), .ZN(new_n230_));
  INV_X1    g029(.A(G92gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(KEYINPUT66), .A3(new_n204_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n227_), .A2(new_n219_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT68), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n226_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n219_), .A2(new_n237_), .A3(new_n224_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(new_n233_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT8), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n239_), .A3(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT67), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n238_), .A2(new_n239_), .A3(new_n246_), .A4(new_n235_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n223_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n236_), .A2(new_n245_), .A3(new_n242_), .A4(new_n247_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(KEYINPUT69), .A3(new_n223_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G57gat), .B(G64gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT11), .ZN(new_n255_));
  XOR2_X1   g054(.A(G71gat), .B(G78gat), .Z(new_n256_));
  OR2_X1    g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n254_), .A2(KEYINPUT11), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n251_), .A2(new_n253_), .A3(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n252_), .A2(new_n223_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n261_), .B1(new_n265_), .B2(new_n260_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n252_), .A2(new_n223_), .A3(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n268_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n265_), .A2(new_n260_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n267_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G120gat), .B(G148gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n275_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT13), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n281_), .B(KEYINPUT13), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT71), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G29gat), .B(G36gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G43gat), .B(G50gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(KEYINPUT76), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(KEYINPUT76), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  OR3_X1    g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n292_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G229gat), .A2(G233gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n292_), .A2(new_n302_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n290_), .B(KEYINPUT15), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n302_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n307_), .A2(new_n304_), .A3(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G113gat), .B(G141gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT82), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G169gat), .B(G197gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n306_), .B2(new_n310_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n285_), .A2(new_n287_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(G197gat), .B(G204gat), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT21), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  OR3_X1    g128(.A1(new_n325_), .A2(new_n328_), .A3(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G228gat), .A2(G233gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT91), .Z(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(KEYINPUT92), .B2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G155gat), .B(G162gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT89), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n337_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(KEYINPUT2), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G141gat), .ZN(new_n341_));
  INV_X1    g140(.A(G148gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n343_), .A2(KEYINPUT3), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(KEYINPUT3), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n344_), .B(new_n345_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n336_), .B1(new_n340_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(KEYINPUT1), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n349_), .B2(KEYINPUT1), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n349_), .A2(new_n352_), .A3(KEYINPUT1), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n343_), .B(new_n348_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n347_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n334_), .B1(new_n357_), .B2(KEYINPUT29), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n333_), .A2(KEYINPUT92), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n347_), .B2(new_n356_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n331_), .ZN(new_n363_));
  OAI211_X1 g162(.A(KEYINPUT92), .B(new_n333_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n322_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n322_), .A3(new_n364_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT90), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n357_), .B2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n347_), .A2(new_n371_), .A3(new_n361_), .A4(new_n356_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G22gat), .B(G50gat), .Z(new_n375_));
  NAND3_X1  g174(.A1(new_n370_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n375_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n368_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n365_), .A2(KEYINPUT94), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  AOI211_X1 g180(.A(new_n381_), .B(new_n322_), .C1(new_n360_), .C2(new_n364_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n367_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n377_), .A2(new_n378_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(KEYINPUT93), .A2(new_n379_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n368_), .B(new_n387_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390_));
  NOR2_X1   g189(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G169gat), .ZN(new_n392_));
  INV_X1    g191(.A(G183gat), .ZN(new_n393_));
  INV_X1    g192(.A(G190gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT23), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(KEYINPUT83), .B(KEYINPUT23), .C1(new_n393_), .C2(new_n394_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G183gat), .A3(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n392_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n395_), .B(KEYINPUT84), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n401_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(G169gat), .B2(G176gat), .ZN(new_n409_));
  NOR3_X1   g208(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT26), .B(G190gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT25), .B(G183gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT95), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n407_), .B(new_n411_), .C1(new_n413_), .C2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n405_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n331_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n407_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n392_), .B1(new_n419_), .B2(new_n404_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n412_), .A2(new_n414_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n402_), .A2(new_n411_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n418_), .B(KEYINPUT20), .C1(new_n331_), .C2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT19), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n423_), .B2(new_n331_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n405_), .A2(new_n416_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(new_n363_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n424_), .A2(new_n426_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT18), .ZN(new_n433_));
  XOR2_X1   g232(.A(G64gat), .B(G92gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n431_), .A2(new_n435_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n390_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n435_), .B(KEYINPUT102), .Z(new_n439_));
  INV_X1    g238(.A(new_n426_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT101), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n331_), .B1(new_n417_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(new_n441_), .B2(new_n417_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n440_), .B1(new_n443_), .B2(new_n428_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n424_), .A2(new_n426_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n439_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n431_), .A2(new_n435_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(KEYINPUT27), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n438_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n389_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G127gat), .B(G134gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT85), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G120gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n357_), .A2(new_n454_), .ZN(new_n455_));
  OR3_X1    g254(.A1(new_n455_), .A2(KEYINPUT97), .A3(KEYINPUT4), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n357_), .A2(new_n454_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(KEYINPUT4), .A3(new_n455_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT96), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT97), .B1(new_n455_), .B2(KEYINPUT4), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n456_), .A2(new_n458_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n457_), .A2(new_n455_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n459_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT99), .ZN(new_n467_));
  XOR2_X1   g266(.A(G57gat), .B(G85gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n465_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n462_), .A2(new_n464_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G71gat), .B(G99gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G43gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n423_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G227gat), .A2(G233gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n480_), .B(G15gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT30), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n482_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n454_), .B(KEYINPUT31), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n485_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n479_), .A2(new_n482_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT86), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n450_), .A2(new_n476_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n449_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n443_), .A2(new_n428_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n426_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n445_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n435_), .A2(KEYINPUT32), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n431_), .A2(KEYINPUT100), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT100), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n501_), .B1(new_n431_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n475_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n436_), .A2(new_n437_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n474_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n462_), .A2(KEYINPUT33), .A3(new_n464_), .A4(new_n471_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n471_), .B1(new_n463_), .B2(new_n460_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .A4(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n379_), .A2(KEYINPUT93), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n384_), .A2(new_n385_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n388_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n496_), .A2(new_n476_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n495_), .B1(new_n520_), .B2(new_n494_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n252_), .A2(new_n223_), .A3(new_n290_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT34), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n522_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n252_), .A2(KEYINPUT69), .A3(new_n223_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT69), .B1(new_n252_), .B2(new_n223_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT72), .B1(new_n533_), .B2(new_n308_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n251_), .A2(KEYINPUT72), .A3(new_n253_), .A4(new_n308_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n530_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n525_), .A2(new_n526_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(KEYINPUT36), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n251_), .A2(new_n253_), .A3(new_n308_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n535_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n538_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n522_), .A2(new_n549_), .A3(new_n527_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n544_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  AOI211_X1 g351(.A(KEYINPUT74), .B(new_n550_), .C1(new_n547_), .C2(new_n535_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n539_), .B(new_n543_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n549_), .B1(new_n548_), .B2(new_n530_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n551_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT74), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n548_), .A2(new_n544_), .A3(new_n551_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n542_), .B(KEYINPUT36), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n554_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT75), .B1(new_n559_), .B2(new_n560_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(KEYINPUT37), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564_));
  OAI221_X1 g363(.A(new_n554_), .B1(KEYINPUT75), .B2(new_n564_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n302_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(new_n260_), .Z(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT79), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n575_), .A2(KEYINPUT77), .A3(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n575_), .A2(new_n576_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n569_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n569_), .A2(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT80), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n321_), .A2(new_n521_), .A3(new_n566_), .A4(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT103), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n475_), .A2(KEYINPUT104), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n475_), .A2(KEYINPUT104), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n294_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT38), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n516_), .A2(new_n519_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n449_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n389_), .A2(new_n476_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n494_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  NOR4_X1   g394(.A1(new_n389_), .A2(new_n493_), .A3(new_n475_), .A4(new_n449_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n561_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n581_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n285_), .A2(new_n287_), .A3(new_n599_), .A4(new_n319_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n476_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n589_), .A2(new_n590_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n591_), .A2(new_n603_), .A3(new_n604_), .ZN(G1324gat));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n601_), .A3(new_n449_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT106), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n607_), .A3(G8gat), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n597_), .A2(new_n593_), .A3(new_n600_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT106), .B1(new_n609_), .B2(new_n295_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n610_), .A3(KEYINPUT39), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT106), .B(new_n612_), .C1(new_n609_), .C2(new_n295_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT105), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n593_), .A2(G8gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n585_), .B2(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n585_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n614_), .B(KEYINPUT40), .C1(new_n617_), .C2(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1325gat));
  OAI21_X1  g422(.A(G15gat), .B1(new_n602_), .B2(new_n493_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT41), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n584_), .A2(G15gat), .A3(new_n493_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1326gat));
  OAI21_X1  g426(.A(G22gat), .B1(new_n602_), .B2(new_n519_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT42), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n519_), .A2(G22gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n584_), .B2(new_n630_), .ZN(G1327gat));
  NAND2_X1  g430(.A1(new_n592_), .A2(new_n594_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n596_), .B1(new_n632_), .B2(new_n493_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n561_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n582_), .A2(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n633_), .A2(new_n320_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n475_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n563_), .A2(new_n565_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n521_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n583_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n521_), .A2(KEYINPUT43), .A3(new_n638_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n321_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n641_), .A2(KEYINPUT44), .A3(new_n321_), .A4(new_n642_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n588_), .A2(G29gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n637_), .B1(new_n647_), .B2(new_n648_), .ZN(G1328gat));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n449_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(G36gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n636_), .A2(new_n652_), .A3(new_n449_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT45), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n651_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  AOI21_X1  g459(.A(G43gat), .B1(new_n636_), .B2(new_n494_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT108), .Z(new_n662_));
  NAND4_X1  g461(.A1(new_n645_), .A2(G43gat), .A3(new_n494_), .A4(new_n646_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g464(.A(G50gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n636_), .A2(new_n666_), .A3(new_n389_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n645_), .A2(new_n389_), .A3(new_n646_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT109), .B1(new_n668_), .B2(G50gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(G1331gat));
  NAND2_X1  g470(.A1(new_n285_), .A2(new_n287_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n319_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n675_), .A2(new_n582_), .A3(new_n597_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(G57gat), .A3(new_n475_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT111), .Z(new_n678_));
  NOR4_X1   g477(.A1(new_n675_), .A2(new_n633_), .A3(new_n638_), .A4(new_n582_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n588_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT110), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT110), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n678_), .A2(new_n681_), .A3(new_n682_), .ZN(G1332gat));
  INV_X1    g482(.A(G64gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n676_), .B2(new_n449_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n679_), .A2(new_n684_), .A3(new_n449_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1333gat));
  INV_X1    g488(.A(G71gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n676_), .B2(new_n494_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT49), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n679_), .A2(new_n690_), .A3(new_n494_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1334gat));
  INV_X1    g493(.A(G78gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n676_), .B2(new_n389_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT50), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n389_), .A2(new_n695_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT113), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n679_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1335gat));
  NOR3_X1   g500(.A1(new_n675_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G85gat), .B1(new_n702_), .B2(new_n588_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT114), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n641_), .A2(new_n642_), .A3(new_n674_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n705_), .A2(new_n230_), .A3(new_n476_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1336gat));
  OAI21_X1  g506(.A(G92gat), .B1(new_n705_), .B2(new_n593_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n231_), .A3(new_n449_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1337gat));
  NAND3_X1  g509(.A1(new_n702_), .A2(new_n220_), .A3(new_n494_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n641_), .A2(new_n494_), .A3(new_n642_), .A4(new_n674_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n712_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT115), .B1(new_n712_), .B2(G99gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g515(.A1(new_n702_), .A2(new_n221_), .A3(new_n389_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n641_), .A2(new_n389_), .A3(new_n642_), .A4(new_n674_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G106gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G106gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g522(.A1(new_n307_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n316_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n311_), .A2(new_n316_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n281_), .A2(new_n726_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n275_), .A2(new_n280_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n319_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n271_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n270_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n264_), .A2(new_n266_), .A3(KEYINPUT55), .A4(new_n269_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n280_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n729_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT116), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n727_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n729_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n739_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT56), .B1(new_n735_), .B2(new_n280_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n743_), .B(new_n741_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n561_), .B1(new_n742_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT57), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n749_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n728_), .A2(new_n726_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n739_), .B1(new_n745_), .B2(KEYINPUT117), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n754_), .B(KEYINPUT56), .C1(new_n735_), .C2(new_n280_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT58), .B(new_n752_), .C1(new_n753_), .C2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT118), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n738_), .A2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n745_), .A2(KEYINPUT117), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n739_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(KEYINPUT58), .A4(new_n752_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n752_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n638_), .A2(new_n757_), .A3(new_n762_), .A4(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n750_), .A2(new_n751_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n319_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n566_), .A2(new_n583_), .A3(new_n768_), .A4(new_n286_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT54), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n769_), .A2(KEYINPUT54), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n767_), .A2(new_n581_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n450_), .A2(new_n494_), .A3(new_n588_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT59), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n748_), .A2(new_n749_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n766_), .A2(new_n751_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n766_), .A2(new_n751_), .A3(KEYINPUT119), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n583_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n771_), .A2(new_n770_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n773_), .A2(KEYINPUT59), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n774_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G113gat), .B1(new_n785_), .B2(new_n768_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n772_), .A2(new_n773_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n319_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1340gat));
  OAI21_X1  g589(.A(G120gat), .B1(new_n785_), .B2(new_n673_), .ZN(new_n791_));
  INV_X1    g590(.A(G120gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n673_), .B2(KEYINPUT60), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n787_), .B(new_n793_), .C1(KEYINPUT60), .C2(new_n792_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(G1341gat));
  NOR3_X1   g594(.A1(new_n772_), .A2(new_n582_), .A3(new_n773_), .ZN(new_n796_));
  OR3_X1    g595(.A1(new_n796_), .A2(KEYINPUT120), .A3(G127gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT120), .B1(new_n796_), .B2(G127gat), .ZN(new_n798_));
  INV_X1    g597(.A(G127gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT121), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n799_), .A2(KEYINPUT121), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n581_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n774_), .B(new_n802_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n797_), .A2(new_n798_), .A3(new_n803_), .ZN(G1342gat));
  OAI21_X1  g603(.A(G134gat), .B1(new_n785_), .B2(new_n566_), .ZN(new_n805_));
  INV_X1    g604(.A(G134gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n787_), .A2(new_n806_), .A3(new_n634_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1343gat));
  NAND2_X1  g607(.A1(new_n767_), .A2(new_n581_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n781_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n496_), .A2(new_n588_), .A3(new_n493_), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(KEYINPUT122), .Z(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n319_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT123), .B(G141gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1344gat));
  NOR2_X1   g616(.A1(new_n813_), .A2(new_n673_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(new_n342_), .ZN(G1345gat));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n583_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT61), .B(G155gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1346gat));
  INV_X1    g621(.A(G162gat), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n813_), .A2(new_n823_), .A3(new_n566_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n813_), .B2(new_n561_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT124), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n827_), .B(new_n823_), .C1(new_n813_), .C2(new_n561_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n824_), .B1(new_n826_), .B2(new_n828_), .ZN(G1347gat));
  INV_X1    g628(.A(KEYINPUT22), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n588_), .A2(new_n593_), .A3(new_n493_), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT125), .Z(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n389_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n319_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n830_), .B(new_n835_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n836_));
  INV_X1    g635(.A(G169gat), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(KEYINPUT62), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(KEYINPUT62), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n778_), .A2(new_n779_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n582_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n834_), .B1(new_n841_), .B2(new_n781_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n837_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n838_), .B1(new_n839_), .B2(new_n844_), .ZN(G1348gat));
  INV_X1    g644(.A(new_n833_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n783_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n672_), .ZN(new_n848_));
  INV_X1    g647(.A(G176gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n772_), .A2(new_n389_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n832_), .A2(new_n849_), .A3(new_n673_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n848_), .A2(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1349gat));
  NOR2_X1   g651(.A1(new_n832_), .A2(new_n582_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G183gat), .B1(new_n850_), .B2(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n599_), .A2(new_n415_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n847_), .B2(new_n855_), .ZN(G1350gat));
  NAND3_X1  g655(.A1(new_n847_), .A2(new_n634_), .A3(new_n412_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n783_), .A2(new_n566_), .A3(new_n846_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n394_), .B2(new_n858_), .ZN(G1351gat));
  NOR4_X1   g658(.A1(new_n494_), .A2(new_n519_), .A3(new_n593_), .A4(new_n475_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n810_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n319_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g663(.A1(new_n861_), .A2(new_n673_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1353gat));
  AOI21_X1  g666(.A(new_n581_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT127), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n869_), .B(new_n872_), .ZN(G1354gat));
  OR3_X1    g672(.A1(new_n861_), .A2(G218gat), .A3(new_n561_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G218gat), .B1(new_n861_), .B2(new_n566_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1355gat));
endmodule


