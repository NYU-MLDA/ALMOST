//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202_));
  INV_X1    g001(.A(G50gat), .ZN(new_n203_));
  INV_X1    g002(.A(G29gat), .ZN(new_n204_));
  INV_X1    g003(.A(G36gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G43gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n207_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n203_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT70), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G43gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G50gat), .A3(new_n209_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n213_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n202_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(new_n216_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT70), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT15), .A3(new_n217_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G1gat), .ZN(new_n225_));
  INV_X1    g024(.A(G8gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT14), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G15gat), .ZN(new_n228_));
  INV_X1    g027(.A(G22gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G15gat), .A2(G22gat), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n227_), .A2(KEYINPUT74), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(KEYINPUT74), .B2(new_n227_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G1gat), .B(G8gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT75), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n233_), .B(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n224_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n221_), .B(KEYINPUT77), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n238_), .B(new_n236_), .Z(new_n242_));
  OAI21_X1  g041(.A(new_n241_), .B1(new_n242_), .B2(new_n240_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244_));
  INV_X1    g043(.A(G169gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G197gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n241_), .B(new_n250_), .C1(new_n242_), .C2(new_n240_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT23), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n257_), .B(new_n259_), .C1(G183gat), .C2(G190gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT22), .B1(new_n262_), .B2(new_n245_), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT22), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT80), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n263_), .A2(new_n269_), .A3(new_n264_), .A4(new_n266_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n260_), .A2(new_n261_), .A3(new_n268_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n245_), .A2(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n261_), .ZN(new_n273_));
  MUX2_X1   g072(.A(new_n272_), .B(new_n273_), .S(KEYINPUT24), .Z(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n253_), .A2(KEYINPUT23), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n255_), .A2(new_n256_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(KEYINPUT23), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n274_), .A2(new_n277_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n271_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G43gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(G127gat), .B(G134gat), .Z(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT83), .B(G113gat), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G120gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT83), .B(G113gat), .ZN(new_n289_));
  INV_X1    g088(.A(G120gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT31), .Z(new_n296_));
  AOI21_X1  g095(.A(new_n285_), .B1(new_n296_), .B2(KEYINPUT82), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(KEYINPUT82), .A3(new_n285_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n284_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n299_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n284_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n302_), .A2(new_n297_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G71gat), .B(G99gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315_));
  INV_X1    g114(.A(new_n294_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT93), .B1(new_n316_), .B2(new_n292_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT93), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n293_), .A2(new_n318_), .A3(new_n294_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(KEYINPUT86), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(KEYINPUT86), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G141gat), .ZN(new_n328_));
  INV_X1    g127(.A(G148gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT3), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(G141gat), .B2(G148gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n323_), .A2(KEYINPUT86), .A3(new_n324_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT87), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n327_), .A2(new_n333_), .A3(new_n337_), .A4(new_n334_), .ZN(new_n338_));
  AOI211_X1 g137(.A(new_n321_), .B(new_n322_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT84), .B1(new_n320_), .B2(KEYINPUT1), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n340_), .A2(new_n322_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n320_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n320_), .B2(KEYINPUT1), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n320_), .A2(new_n343_), .A3(KEYINPUT1), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n328_), .A2(new_n329_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n323_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n317_), .B(new_n319_), .C1(new_n339_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n336_), .A2(new_n338_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n322_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n320_), .A3(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n353_), .A2(KEYINPUT93), .A3(new_n295_), .A4(new_n348_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n315_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n322_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n349_), .B1(new_n356_), .B2(new_n320_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n295_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n357_), .A2(KEYINPUT4), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n314_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n350_), .A2(new_n313_), .A3(new_n354_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G1gat), .B(G29gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n360_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n312_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n353_), .A2(new_n348_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G22gat), .B(G50gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT28), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n374_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G228gat), .ZN(new_n378_));
  INV_X1    g177(.A(G233gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n247_), .A2(G204gat), .ZN(new_n383_));
  INV_X1    g182(.A(G204gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(G197gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT21), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(G197gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n247_), .A2(G204gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT21), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G211gat), .A2(G218gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G211gat), .A2(G218gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT88), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(G211gat), .A2(G218gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n391_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n386_), .A2(new_n390_), .A3(new_n394_), .A4(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n389_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n392_), .A2(new_n393_), .A3(KEYINPUT88), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n395_), .B2(new_n391_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT89), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n402_), .A3(KEYINPUT89), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n381_), .B1(new_n382_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT90), .Z(new_n410_));
  NAND2_X1  g209(.A1(new_n403_), .A2(new_n381_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n373_), .B2(KEYINPUT29), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n408_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n410_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n412_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n353_), .B2(new_n348_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n407_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n380_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n414_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n377_), .B1(new_n413_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n409_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n407_), .B1(new_n357_), .B2(new_n416_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n412_), .B1(new_n423_), .B2(new_n380_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n422_), .A2(KEYINPUT91), .B1(new_n414_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n374_), .B(new_n376_), .Z(new_n426_));
  NAND4_X1  g225(.A1(new_n415_), .A2(new_n419_), .A3(KEYINPUT91), .A4(new_n414_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n421_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT92), .Z(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT19), .Z(new_n433_));
  NAND4_X1  g232(.A1(new_n274_), .A2(new_n277_), .A3(new_n259_), .A4(new_n257_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT22), .B(G169gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n264_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n278_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n256_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n440_), .B2(new_n258_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G183gat), .A2(G190gat), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n261_), .B(new_n436_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n405_), .A2(new_n406_), .A3(new_n434_), .A4(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n282_), .A2(new_n403_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT95), .B1(new_n444_), .B2(KEYINPUT20), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n433_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n434_), .A2(new_n443_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n403_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n433_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n403_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n281_), .A3(new_n271_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n451_), .A2(KEYINPUT20), .A3(new_n452_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT18), .B(G64gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G92gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(new_n434_), .A3(new_n443_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n446_), .A2(new_n462_), .A3(KEYINPUT20), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n452_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n451_), .A2(KEYINPUT20), .A3(new_n433_), .A4(new_n454_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n460_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n461_), .A2(KEYINPUT27), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n372_), .A2(new_n430_), .A3(new_n474_), .ZN(new_n475_));
  AND4_X1   g274(.A1(new_n370_), .A2(new_n429_), .A3(new_n473_), .A4(new_n469_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n456_), .B2(new_n477_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT96), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT96), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n479_), .B(new_n482_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n360_), .A2(new_n361_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n366_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n350_), .A2(new_n354_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n366_), .B1(new_n488_), .B2(new_n314_), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n355_), .A2(new_n314_), .A3(new_n359_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n471_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n369_), .A2(KEYINPUT33), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n481_), .A2(new_n483_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n476_), .B1(new_n494_), .B2(new_n430_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n312_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n475_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT10), .B(G99gat), .Z(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(KEYINPUT9), .A3(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT6), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n500_), .A2(new_n503_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n508_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513_));
  INV_X1    g312(.A(G99gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n499_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(KEYINPUT65), .A3(new_n509_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n506_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n501_), .A2(new_n502_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT64), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT64), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n501_), .A2(new_n520_), .A3(new_n502_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n517_), .A2(KEYINPUT66), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT66), .B1(new_n517_), .B2(new_n522_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n506_), .A2(new_n515_), .A3(new_n509_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n221_), .B(new_n507_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n220_), .A2(new_n223_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n507_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n517_), .A2(new_n522_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT66), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n517_), .A2(KEYINPUT66), .A3(new_n522_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(KEYINPUT8), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n532_), .B1(new_n537_), .B2(new_n528_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n530_), .B1(new_n531_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT34), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n539_), .A2(KEYINPUT71), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n539_), .B2(KEYINPUT71), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n542_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT72), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n537_), .A2(new_n528_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n550_), .A2(new_n507_), .B1(new_n223_), .B2(new_n220_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n221_), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n532_), .B(new_n552_), .C1(new_n537_), .C2(new_n528_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT71), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n544_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n539_), .A2(KEYINPUT71), .A3(new_n545_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(KEYINPUT35), .A3(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n548_), .A2(new_n549_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G134gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G162gat), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n548_), .A2(new_n549_), .A3(new_n557_), .A4(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n546_), .A2(new_n547_), .A3(new_n540_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n541_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n567_));
  OAI211_X1 g366(.A(KEYINPUT36), .B(new_n561_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT73), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n507_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G57gat), .B(G64gat), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT11), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT11), .ZN(new_n576_));
  XOR2_X1   g375(.A(G71gat), .B(G78gat), .Z(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n576_), .A2(new_n577_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n550_), .A2(new_n507_), .A3(new_n580_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT67), .A3(new_n583_), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n573_), .A2(KEYINPUT67), .A3(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  AOI211_X1 g387(.A(new_n532_), .B(new_n581_), .C1(new_n537_), .C2(new_n528_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT68), .B1(new_n589_), .B2(new_n587_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n591_), .B1(new_n538_), .B2(new_n580_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT68), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n583_), .A2(new_n593_), .A3(new_n586_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n573_), .A2(KEYINPUT12), .A3(new_n581_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(new_n592_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n588_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G120gat), .B(G148gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n597_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(KEYINPUT13), .A3(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n580_), .B(new_n613_), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n236_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT16), .B(G183gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  NOR3_X1   g419(.A1(new_n615_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(KEYINPUT17), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n615_), .B2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n569_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n572_), .A2(new_n612_), .A3(new_n623_), .A4(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT76), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n252_), .B(new_n497_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n626_), .B2(new_n625_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n225_), .A3(new_n371_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT97), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n569_), .B(KEYINPUT98), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n635_), .A2(new_n497_), .A3(new_n623_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n252_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n611_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(new_n371_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n632_), .B(new_n633_), .C1(new_n225_), .C2(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n474_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n226_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT39), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n628_), .A2(new_n226_), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g446(.A(new_n228_), .B1(new_n639_), .B2(new_n496_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n628_), .A2(new_n228_), .A3(new_n496_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  OR2_X1    g450(.A1(new_n430_), .A2(KEYINPUT99), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n430_), .A2(KEYINPUT99), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n229_), .B1(new_n639_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT42), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n628_), .A2(new_n229_), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1327gat));
  AND2_X1   g458(.A1(new_n497_), .A2(new_n569_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n611_), .A2(new_n637_), .A3(new_n623_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n204_), .A3(new_n371_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n572_), .A2(new_n624_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n497_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n497_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n624_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT37), .B1(new_n569_), .B2(KEYINPUT73), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT101), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n572_), .A2(new_n674_), .A3(new_n624_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT100), .B(new_n475_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n670_), .A2(new_n673_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT102), .B1(new_n677_), .B2(KEYINPUT43), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n668_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n665_), .B1(new_n680_), .B2(new_n661_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n683_), .A3(new_n661_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n370_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n663_), .B1(new_n685_), .B2(new_n204_), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n680_), .A2(new_n661_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n688_), .B2(new_n665_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n205_), .B1(new_n689_), .B2(new_n642_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n662_), .A2(new_n205_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(KEYINPUT104), .A3(new_n474_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT104), .B1(new_n691_), .B2(new_n474_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(KEYINPUT45), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT45), .B1(new_n693_), .B2(new_n694_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n687_), .B1(new_n690_), .B2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n695_), .A2(new_n696_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n474_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n699_), .B(KEYINPUT46), .C1(new_n700_), .C2(new_n205_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1329gat));
  XNOR2_X1  g501(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT106), .Z(new_n704_));
  AND3_X1   g503(.A1(new_n680_), .A2(new_n683_), .A3(new_n661_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n496_), .B1(new_n705_), .B2(new_n681_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G43gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n662_), .A2(new_n207_), .A3(new_n496_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n704_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n708_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n710_), .B(new_n711_), .C1(new_n706_), .C2(G43gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1330gat));
  NAND2_X1  g512(.A1(new_n655_), .A2(new_n203_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n662_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n430_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n203_), .ZN(G1331gat));
  INV_X1    g517(.A(new_n623_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n671_), .A2(new_n672_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n611_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n637_), .B(new_n497_), .C1(new_n721_), .C2(KEYINPUT108), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(KEYINPUT108), .B2(new_n721_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n371_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT109), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n612_), .A2(new_n252_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n636_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n371_), .A2(G57gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1332gat));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n642_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G64gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT110), .Z(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT48), .ZN(new_n733_));
  INV_X1    g532(.A(new_n723_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n734_), .A2(G64gat), .A3(new_n474_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n727_), .B2(new_n496_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT49), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n723_), .A2(new_n737_), .A3(new_n496_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1334gat));
  NAND2_X1  g540(.A1(new_n727_), .A2(new_n655_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G78gat), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT111), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT50), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n654_), .A2(G78gat), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT112), .Z(new_n747_));
  OAI21_X1  g546(.A(new_n745_), .B1(new_n734_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n726_), .A2(new_n719_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n660_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT113), .Z(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n371_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT114), .Z(new_n754_));
  AND2_X1   g553(.A1(new_n680_), .A2(new_n750_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n371_), .A2(G85gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  AOI21_X1  g556(.A(G92gat), .B1(new_n752_), .B2(new_n642_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n642_), .A2(G92gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n755_), .B2(new_n759_), .ZN(G1337gat));
  AOI21_X1  g559(.A(new_n514_), .B1(new_n755_), .B2(new_n496_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n752_), .A2(new_n498_), .A3(new_n496_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n752_), .A2(new_n499_), .A3(new_n429_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n680_), .A2(new_n429_), .A3(new_n750_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n767_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n720_), .A2(new_n777_), .A3(new_n637_), .A4(new_n612_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT54), .B1(new_n625_), .B2(new_n252_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n595_), .A2(new_n592_), .A3(new_n583_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT115), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n595_), .A2(new_n592_), .A3(new_n783_), .A4(new_n583_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n587_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n596_), .A2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n595_), .A2(new_n592_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(KEYINPUT55), .A3(new_n590_), .A4(new_n594_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n603_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(new_n240_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n237_), .A2(new_n793_), .A3(new_n239_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n248_), .C1(new_n242_), .C2(new_n793_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(new_n251_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n790_), .A2(new_n797_), .A3(new_n603_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n792_), .A2(new_n605_), .A3(new_n796_), .A4(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT117), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT58), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT117), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n666_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n791_), .A2(KEYINPUT116), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n790_), .A2(new_n806_), .A3(new_n797_), .A4(new_n603_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n637_), .A2(new_n604_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n792_), .A2(new_n805_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n607_), .A2(new_n796_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n569_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n804_), .A2(new_n815_), .A3(KEYINPUT119), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT119), .B1(new_n804_), .B2(new_n815_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n812_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n816_), .A2(new_n817_), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n780_), .B1(new_n820_), .B2(new_n623_), .ZN(new_n821_));
  NOR4_X1   g620(.A1(new_n642_), .A2(new_n312_), .A3(new_n370_), .A4(new_n429_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n812_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n798_), .A2(new_n796_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n604_), .B1(new_n791_), .B2(KEYINPUT56), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n827_), .B(KEYINPUT58), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n802_), .B1(new_n799_), .B2(KEYINPUT117), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n826_), .B1(new_n832_), .B2(new_n666_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n623_), .B1(new_n833_), .B2(new_n818_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n778_), .A2(new_n779_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT118), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n804_), .A2(new_n815_), .A3(new_n818_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n719_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n780_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n840_), .A3(new_n822_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n825_), .B(new_n252_), .C1(new_n842_), .C2(new_n823_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G113gat), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n841_), .A2(G113gat), .A3(new_n637_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n845_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n841_), .A2(KEYINPUT59), .B1(new_n821_), .B2(new_n824_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n252_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT120), .B1(new_n851_), .B2(new_n846_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n852_), .ZN(G1340gat));
  OAI211_X1 g652(.A(new_n825_), .B(new_n611_), .C1(new_n842_), .C2(new_n823_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n856_));
  AOI21_X1  g655(.A(G120gat), .B1(new_n611_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n842_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n290_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n855_), .A2(KEYINPUT121), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n290_), .B1(new_n850_), .B2(new_n611_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n857_), .B(new_n841_), .C1(new_n856_), .C2(G120gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n864_), .ZN(G1341gat));
  AOI21_X1  g664(.A(G127gat), .B1(new_n842_), .B2(new_n623_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n850_), .A2(G127gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n623_), .ZN(G1342gat));
  AOI21_X1  g667(.A(G134gat), .B1(new_n842_), .B2(new_n634_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n666_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT122), .B(G134gat), .Z(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n850_), .B2(new_n872_), .ZN(G1343gat));
  NAND4_X1  g672(.A1(new_n836_), .A2(new_n429_), .A3(new_n312_), .A4(new_n840_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n642_), .A2(new_n370_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n252_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n611_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n623_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  NOR3_X1   g683(.A1(new_n874_), .A2(new_n635_), .A3(new_n876_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n838_), .A2(new_n839_), .A3(new_n780_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n839_), .B1(new_n838_), .B2(new_n780_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n496_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(new_n429_), .A3(new_n875_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n673_), .A2(new_n675_), .A3(G162gat), .ZN(new_n890_));
  OAI22_X1  g689(.A1(new_n885_), .A2(G162gat), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT123), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  OAI221_X1 g692(.A(new_n893_), .B1(new_n889_), .B2(new_n890_), .C1(G162gat), .C2(new_n885_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1347gat));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n372_), .A2(new_n642_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n821_), .A2(new_n654_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n252_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n896_), .B1(new_n900_), .B2(G169gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n821_), .A2(new_n654_), .A3(new_n898_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n896_), .B(G169gat), .C1(new_n902_), .C2(new_n637_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n252_), .A2(new_n435_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT124), .Z(new_n906_));
  OAI22_X1  g705(.A1(new_n901_), .A2(new_n904_), .B1(new_n902_), .B2(new_n906_), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n899_), .B2(new_n611_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n886_), .A2(new_n887_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT125), .B1(new_n909_), .B2(new_n430_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n886_), .A2(new_n887_), .A3(new_n911_), .A4(new_n429_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G176gat), .B1(new_n910_), .B2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n612_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n908_), .B1(new_n914_), .B2(new_n898_), .ZN(G1349gat));
  NOR3_X1   g714(.A1(new_n902_), .A2(new_n275_), .A3(new_n719_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n623_), .B(new_n898_), .C1(new_n910_), .C2(new_n912_), .ZN(new_n917_));
  INV_X1    g716(.A(G183gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n899_), .A2(new_n276_), .A3(new_n634_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G190gat), .B1(new_n902_), .B2(new_n870_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT126), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n920_), .A2(new_n924_), .A3(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n430_), .A2(new_n371_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n888_), .A2(KEYINPUT127), .A3(new_n927_), .A4(new_n642_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n836_), .A2(new_n927_), .A3(new_n312_), .A4(new_n840_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n474_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n928_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n252_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G197gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1352gat));
  AOI21_X1  g735(.A(G204gat), .B1(new_n932_), .B2(new_n611_), .ZN(new_n937_));
  AOI211_X1 g736(.A(new_n384_), .B(new_n612_), .C1(new_n928_), .C2(new_n931_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1353gat));
  OR2_X1    g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n940_), .B1(new_n932_), .B2(new_n623_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT63), .B(G211gat), .ZN(new_n942_));
  AOI211_X1 g741(.A(new_n719_), .B(new_n942_), .C1(new_n928_), .C2(new_n931_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n932_), .B2(new_n634_), .ZN(new_n945_));
  INV_X1    g744(.A(G218gat), .ZN(new_n946_));
  AOI211_X1 g745(.A(new_n946_), .B(new_n870_), .C1(new_n928_), .C2(new_n931_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1355gat));
endmodule


