//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT82), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(new_n203_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT82), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT84), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(new_n217_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n216_), .A2(new_n229_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n210_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n207_), .A2(new_n204_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n231_), .A2(new_n232_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n226_), .B(new_n235_), .C1(new_n236_), .C2(new_n228_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n237_), .A3(KEYINPUT4), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT98), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT98), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n234_), .A2(new_n237_), .A3(new_n240_), .A4(KEYINPUT4), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT99), .B1(new_n234_), .B2(KEYINPUT4), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n226_), .B1(new_n236_), .B2(new_n228_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT99), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .A4(new_n210_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n239_), .A2(new_n241_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n234_), .A2(new_n237_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G1gat), .B(G29gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G85gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G57gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n259_), .A3(new_n252_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n227_), .A2(new_n233_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(G228gat), .A2(G233gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT87), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G218gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G211gat), .ZN(new_n272_));
  INV_X1    g071(.A(G211gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G218gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n272_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n270_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n273_), .A2(G218gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n271_), .A2(G211gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT88), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n268_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n283_), .A3(KEYINPUT21), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT89), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n270_), .B(new_n286_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n285_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n266_), .A2(new_n267_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n267_), .B1(new_n266_), .B2(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n284_), .A2(new_n287_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n265_), .B1(new_n264_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT91), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  OAI22_X1  g099(.A1(new_n293_), .A2(new_n294_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G78gat), .B(G106gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G22gat), .B(G50gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT86), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n243_), .B2(KEYINPUT29), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n262_), .A2(new_n263_), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n309_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n302_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n302_), .A2(KEYINPUT92), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n301_), .B(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G71gat), .B(G99gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G43gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT31), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT23), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT77), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G190gat), .ZN(new_n332_));
  INV_X1    g131(.A(G183gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n325_), .A2(KEYINPUT80), .A3(G183gat), .A4(G190gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338_));
  AOI21_X1  g137(.A(G176gat), .B1(new_n338_), .B2(G169gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n340_));
  INV_X1    g139(.A(G169gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n338_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n339_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n343_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n345_), .B(KEYINPUT22), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n336_), .B(new_n337_), .C1(new_n346_), .C2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT24), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n337_), .A2(KEYINPUT24), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n352_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n324_), .A2(new_n326_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT25), .B(G183gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n351_), .A2(KEYINPUT81), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT81), .B1(new_n351_), .B2(new_n364_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(G15gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n351_), .A2(new_n364_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n351_), .A2(KEYINPUT81), .A3(new_n364_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n371_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n210_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n210_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n322_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n321_), .A3(new_n381_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n318_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(G190gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n356_), .B1(new_n359_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n335_), .A3(new_n328_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT22), .B(G169gat), .Z(new_n397_));
  NOR2_X1   g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  OAI221_X1 g197(.A(new_n337_), .B1(new_n397_), .B2(G176gat), .C1(new_n357_), .C2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n295_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n367_), .B2(new_n290_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT94), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n401_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n295_), .A2(KEYINPUT89), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n375_), .A2(new_n406_), .A3(new_n376_), .A4(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n404_), .A3(KEYINPUT20), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n393_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n291_), .A2(new_n377_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n296_), .A2(new_n399_), .A3(new_n396_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n393_), .A2(new_n402_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT96), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n411_), .A2(KEYINPUT97), .A3(new_n416_), .A4(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n401_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n408_), .A2(KEYINPUT20), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n426_), .B2(KEYINPUT94), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n392_), .B1(new_n427_), .B2(new_n409_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n428_), .B2(new_n415_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(KEYINPUT94), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n409_), .A3(new_n401_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n415_), .B1(new_n432_), .B2(new_n393_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT97), .B1(new_n433_), .B2(new_n422_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n389_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT104), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n412_), .A2(new_n413_), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n438_));
  OAI21_X1  g237(.A(new_n393_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n432_), .B2(new_n393_), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n422_), .B(KEYINPUT103), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n422_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT27), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n435_), .A2(new_n436_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n436_), .B1(new_n435_), .B2(new_n444_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n261_), .B(new_n388_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n435_), .A2(new_n261_), .A3(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n318_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n384_), .A2(new_n386_), .A3(KEYINPUT83), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT83), .B1(new_n384_), .B2(new_n386_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n430_), .A2(new_n434_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n247_), .A2(new_n248_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n259_), .B1(new_n251_), .B2(new_n249_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n456_), .B1(new_n260_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT101), .ZN(new_n459_));
  INV_X1    g258(.A(new_n252_), .ZN(new_n460_));
  AOI211_X1 g259(.A(new_n257_), .B(new_n460_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n260_), .A2(KEYINPUT101), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n453_), .A2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n258_), .A2(new_n260_), .B1(new_n440_), .B2(new_n468_), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n428_), .A2(new_n415_), .A3(new_n468_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n318_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n452_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n449_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n447_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G1gat), .ZN(new_n475_));
  INV_X1    g274(.A(G8gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT14), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n483_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n479_), .A2(new_n485_), .A3(new_n480_), .A4(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n487_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n490_), .B(KEYINPUT15), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT75), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n487_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n496_), .A2(new_n487_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT75), .B1(new_n487_), .B2(new_n491_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n495_), .B1(new_n493_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G113gat), .B(G141gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(G169gat), .B(G197gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT76), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n502_), .A2(new_n507_), .A3(new_n505_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G85gat), .B(G92gat), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT9), .ZN(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT9), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n515_), .A2(new_n518_), .A3(new_n520_), .A4(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n519_), .B1(new_n527_), .B2(new_n514_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n528_), .B(KEYINPUT8), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT65), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n524_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT64), .B(G71gat), .ZN(new_n536_));
  INV_X1    g335(.A(G78gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n539_), .B(KEYINPUT11), .Z(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n538_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(KEYINPUT12), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(new_n524_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n543_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT66), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT66), .B1(new_n546_), .B2(new_n547_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n544_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n545_), .A2(new_n543_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT67), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n545_), .A2(new_n543_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  INV_X1    g356(.A(new_n554_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n553_), .A2(new_n546_), .ZN(new_n561_));
  OAI22_X1  g360(.A1(new_n552_), .A2(new_n560_), .B1(new_n554_), .B2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G120gat), .B(G148gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n562_), .A2(new_n567_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT13), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT13), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(KEYINPUT69), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n568_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n562_), .A2(new_n567_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n562_), .A2(new_n567_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT13), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n575_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n511_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n474_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT71), .ZN(new_n585_));
  XOR2_X1   g384(.A(G134gat), .B(G162gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT36), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n533_), .A2(new_n490_), .A3(new_n524_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n535_), .B2(new_n496_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n591_), .A2(KEYINPUT70), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n524_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n533_), .A2(KEYINPUT65), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n530_), .A2(new_n531_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n496_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n589_), .B(KEYINPUT70), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n593_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n595_), .A2(new_n597_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT35), .B1(new_n595_), .B2(new_n604_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n605_), .A2(new_n606_), .A3(KEYINPUT72), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT72), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n594_), .B1(new_n591_), .B2(KEYINPUT70), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n603_), .A2(new_n593_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n596_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n595_), .A2(new_n597_), .A3(new_n604_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(KEYINPUT73), .B(new_n588_), .C1(new_n607_), .C2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n605_), .A2(new_n606_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n587_), .A2(KEYINPUT36), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n588_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT72), .B1(new_n605_), .B2(new_n606_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n611_), .A2(new_n608_), .A3(new_n612_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n620_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(KEYINPUT73), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n583_), .B1(new_n619_), .B2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n618_), .B(KEYINPUT37), .C1(new_n620_), .C2(new_n616_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n487_), .B(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(new_n543_), .Z(new_n630_));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT16), .ZN(new_n632_));
  XOR2_X1   g431(.A(G183gat), .B(G211gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n630_), .B1(KEYINPUT17), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT17), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n634_), .B(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n630_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n627_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n582_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n261_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n475_), .A3(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT105), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n619_), .A2(new_n624_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n640_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n582_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n261_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n647_), .A2(new_n648_), .A3(new_n653_), .ZN(G1324gat));
  NOR2_X1   g453(.A1(new_n445_), .A2(new_n446_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n476_), .B1(new_n657_), .B2(KEYINPUT39), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(KEYINPUT106), .A3(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n656_), .B(new_n658_), .C1(new_n657_), .C2(KEYINPUT39), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n642_), .A2(new_n476_), .A3(new_n655_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1325gat));
  NAND3_X1  g465(.A1(new_n642_), .A2(new_n369_), .A3(new_n452_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT107), .Z(new_n668_));
  AOI21_X1  g467(.A(new_n369_), .B1(new_n651_), .B2(new_n452_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT41), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n318_), .B(KEYINPUT108), .Z(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n651_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT42), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n642_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(new_n649_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n640_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n582_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n643_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n474_), .A2(new_n627_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n685_), .A2(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n474_), .A2(new_n627_), .A3(new_n685_), .A4(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n574_), .A2(new_n580_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n510_), .A3(new_n640_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n581_), .A2(KEYINPUT109), .A3(new_n640_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n688_), .A2(new_n689_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n688_), .A2(new_n695_), .A3(KEYINPUT44), .A4(new_n689_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n643_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n683_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(new_n655_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n582_), .A2(new_n680_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n698_), .A2(new_n655_), .A3(new_n699_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n711_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n709_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1329gat));
  INV_X1    g515(.A(new_n387_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n698_), .A2(G43gat), .A3(new_n717_), .A4(new_n699_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT112), .B(G43gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n452_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n681_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n682_), .B2(new_n673_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n318_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n700_), .B2(new_n725_), .ZN(G1331gat));
  AOI211_X1 g525(.A(new_n510_), .B(new_n690_), .C1(new_n447_), .C2(new_n473_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(new_n641_), .ZN(new_n728_));
  INV_X1    g527(.A(G57gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n643_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n727_), .A2(new_n643_), .A3(new_n650_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n728_), .A2(new_n733_), .A3(new_n655_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n727_), .A2(new_n655_), .A3(new_n650_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G64gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G64gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1333gat));
  NOR2_X1   g538(.A1(new_n720_), .A2(G71gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT113), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n728_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n727_), .A2(new_n452_), .A3(new_n650_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G71gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1334gat));
  NAND3_X1  g546(.A1(new_n728_), .A2(new_n537_), .A3(new_n673_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n727_), .A2(new_n650_), .A3(new_n673_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G78gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G78gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1335gat));
  NOR3_X1   g552(.A1(new_n690_), .A2(new_n510_), .A3(new_n679_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n688_), .A2(new_n689_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n261_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n727_), .A2(new_n680_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n521_), .A3(new_n643_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1336gat));
  OAI21_X1  g559(.A(G92gat), .B1(new_n755_), .B2(new_n703_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n522_), .A3(new_n655_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1337gat));
  OAI21_X1  g562(.A(G99gat), .B1(new_n755_), .B2(new_n720_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n516_), .A3(new_n717_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n766_), .B(new_n767_), .Z(G1338gat));
  NAND4_X1  g567(.A1(new_n688_), .A2(new_n318_), .A3(new_n689_), .A4(new_n754_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n517_), .B1(new_n770_), .B2(KEYINPUT52), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(KEYINPUT115), .A3(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n769_), .B(new_n771_), .C1(new_n770_), .C2(KEYINPUT52), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n758_), .A2(new_n517_), .A3(new_n318_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  INV_X1    g578(.A(new_n627_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT116), .B1(new_n511_), .B2(new_n679_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n510_), .A2(new_n640_), .A3(new_n782_), .ZN(new_n783_));
  NOR4_X1   g582(.A1(new_n576_), .A2(new_n781_), .A3(new_n579_), .A4(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n779_), .B1(new_n780_), .B2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n784_), .A2(new_n625_), .A3(new_n779_), .A4(new_n626_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n787_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n501_), .A2(new_n494_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n505_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n570_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n553_), .B(new_n544_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n558_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT118), .ZN(new_n800_));
  INV_X1    g599(.A(new_n560_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n550_), .A2(new_n551_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(KEYINPUT55), .A4(new_n544_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(new_n804_), .A3(new_n558_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n552_), .B2(new_n560_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n800_), .A2(new_n803_), .A3(new_n805_), .A4(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n797_), .B1(new_n808_), .B2(new_n567_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n577_), .A2(new_n510_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n809_), .B2(KEYINPUT56), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n796_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n649_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n808_), .A2(new_n567_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n567_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(KEYINPUT121), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n821_), .A3(new_n817_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n795_), .A2(new_n569_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n820_), .A2(KEYINPUT58), .A3(new_n822_), .A4(new_n823_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n627_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n815_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n813_), .B2(new_n649_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n640_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n791_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n703_), .A2(new_n643_), .A3(new_n388_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n836_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n831_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n796_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n816_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n845_));
  INV_X1    g644(.A(new_n811_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n844_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n678_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(KEYINPUT120), .A3(new_n830_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n843_), .A2(new_n851_), .A3(new_n815_), .A4(new_n828_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n640_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n839_), .B1(new_n853_), .B2(new_n791_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n841_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n511_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n854_), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n858_), .A2(G113gat), .A3(new_n511_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n856_), .B2(new_n690_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n690_), .A2(KEYINPUT60), .ZN(new_n862_));
  MUX2_X1   g661(.A(new_n862_), .B(KEYINPUT60), .S(G120gat), .Z(new_n863_));
  NAND2_X1  g662(.A1(new_n854_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n856_), .B2(new_n640_), .ZN(new_n866_));
  OR3_X1    g665(.A1(new_n858_), .A2(G127gat), .A3(new_n640_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1342gat));
  OAI21_X1  g667(.A(G134gat), .B1(new_n856_), .B2(new_n780_), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n858_), .A2(G134gat), .A3(new_n678_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1343gat));
  AND2_X1   g670(.A1(new_n720_), .A2(new_n318_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n655_), .A2(new_n873_), .A3(new_n261_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n853_), .B2(new_n791_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n510_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n876_), .A2(new_n879_), .A3(new_n510_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT123), .B(G141gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n881_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n876_), .B2(new_n510_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n640_), .A2(new_n852_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n885_));
  NOR4_X1   g684(.A1(new_n885_), .A2(KEYINPUT124), .A3(new_n511_), .A4(new_n875_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n887_), .ZN(G1344gat));
  INV_X1    g687(.A(new_n690_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n876_), .A2(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g690(.A1(new_n876_), .A2(new_n679_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  AOI21_X1  g693(.A(G162gat), .B1(new_n876_), .B2(new_n649_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n627_), .A2(G162gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT125), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n876_), .B2(new_n897_), .ZN(G1347gat));
  NAND2_X1  g697(.A1(new_n655_), .A2(new_n261_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n720_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n673_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n834_), .A2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903_), .B2(new_n511_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(G169gat), .C1(new_n903_), .C2(new_n511_), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n903_), .A2(new_n511_), .A3(new_n397_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1348gat));
  INV_X1    g708(.A(G176gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n834_), .A2(new_n889_), .A3(new_n902_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n885_), .A2(new_n318_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n901_), .A2(new_n910_), .A3(new_n690_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n910_), .A2(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1349gat));
  NOR3_X1   g713(.A1(new_n903_), .A2(new_n359_), .A3(new_n640_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(new_n679_), .A3(new_n900_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n333_), .B2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n903_), .B2(new_n780_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n649_), .A2(new_n394_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n903_), .B2(new_n919_), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n899_), .A2(new_n873_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n885_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n510_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g724(.A1(new_n885_), .A2(new_n690_), .A3(new_n922_), .ZN(new_n926_));
  INV_X1    g725(.A(G204gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(KEYINPUT127), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(KEYINPUT120), .B1(new_n850_), .B2(new_n830_), .ZN(new_n929_));
  AOI211_X1 g728(.A(new_n842_), .B(KEYINPUT57), .C1(new_n849_), .C2(new_n678_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n824_), .A2(new_n825_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n932_));
  AOI22_X1  g731(.A1(new_n827_), .A2(new_n932_), .B1(new_n814_), .B2(KEYINPUT57), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n679_), .B1(new_n931_), .B2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n790_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n935_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n889_), .B(new_n921_), .C1(new_n934_), .C2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n937_), .A2(new_n938_), .A3(G204gat), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n937_), .A2(new_n940_), .A3(G204gat), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n937_), .B2(G204gat), .ZN(new_n942_));
  OAI22_X1  g741(.A1(new_n928_), .A2(new_n939_), .B1(new_n941_), .B2(new_n942_), .ZN(G1353gat));
  OAI21_X1  g742(.A(new_n921_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  AND2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  NOR4_X1   g745(.A1(new_n944_), .A2(new_n640_), .A3(new_n945_), .A4(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n923_), .A2(new_n679_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n945_), .ZN(G1354gat));
  NAND3_X1  g748(.A1(new_n923_), .A2(new_n271_), .A3(new_n649_), .ZN(new_n950_));
  OAI21_X1  g749(.A(G218gat), .B1(new_n944_), .B2(new_n780_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1355gat));
endmodule


