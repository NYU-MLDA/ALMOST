//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  XOR2_X1   g000(.A(G22gat), .B(G50gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OR4_X1    g002(.A1(KEYINPUT83), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n208_));
  OAI22_X1  g007(.A1(KEYINPUT83), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT80), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT81), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(new_n212_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n215_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT82), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(new_n219_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n212_), .B(KEYINPUT82), .C1(new_n215_), .C2(new_n219_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G141gat), .B(G148gat), .Z(new_n226_));
  AOI21_X1  g025(.A(new_n218_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT28), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT28), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n203_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n231_), .A3(new_n203_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n225_), .A2(new_n226_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n217_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT87), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT29), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT85), .ZN(new_n240_));
  INV_X1    g039(.A(G197gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(G204gat), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G211gat), .B(G218gat), .Z(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  OAI221_X1 g043(.A(new_n242_), .B1(new_n241_), .B2(G204gat), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n243_), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n248_));
  AOI211_X1 g047(.A(KEYINPUT86), .B(new_n244_), .C1(G197gat), .C2(G204gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n243_), .B1(KEYINPUT86), .B2(new_n244_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n240_), .A2(new_n241_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n245_), .A2(new_n250_), .A3(new_n251_), .A4(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT87), .B1(new_n227_), .B2(new_n228_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n239_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G228gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n237_), .A2(KEYINPUT84), .A3(KEYINPUT29), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n260_), .A2(new_n262_), .A3(new_n257_), .A4(new_n254_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n259_), .A2(KEYINPUT89), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT89), .B1(new_n259_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n235_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n259_), .A2(KEYINPUT89), .A3(new_n263_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(KEYINPUT88), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n271_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n266_), .A2(new_n273_), .A3(new_n268_), .ZN(new_n274_));
  INV_X1    g073(.A(G120gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G113gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n276_), .A2(G113gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n275_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n276_), .A2(G113gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(G120gat), .A3(new_n277_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n237_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n227_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(KEYINPUT4), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n227_), .A2(KEYINPUT4), .A3(new_n285_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n284_), .A2(new_n288_), .A3(new_n286_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT0), .B(G57gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(G85gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(G1gat), .B(G29gat), .Z(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n292_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  INV_X1    g102(.A(G183gat), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n306_), .B(new_n307_), .C1(G183gat), .C2(G190gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT77), .B(G176gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT22), .B(G169gat), .Z(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n309_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n306_), .A2(new_n307_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT26), .B(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(KEYINPUT76), .A3(G183gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT25), .B1(new_n317_), .B2(new_n304_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G169gat), .ZN(new_n320_));
  INV_X1    g119(.A(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(KEYINPUT24), .A3(new_n309_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(KEYINPUT24), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n313_), .A2(new_n319_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n312_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n312_), .B2(new_n325_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n254_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n314_), .ZN(new_n330_));
  XOR2_X1   g129(.A(KEYINPUT25), .B(G183gat), .Z(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n332_), .A2(new_n323_), .A3(new_n324_), .A4(new_n313_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n311_), .A2(new_n310_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n309_), .A2(KEYINPUT91), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n309_), .A2(KEYINPUT91), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n308_), .A4(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n253_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n329_), .A2(KEYINPUT20), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT90), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT19), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n328_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n312_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n253_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n333_), .A2(new_n337_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n254_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(KEYINPUT20), .A3(new_n342_), .A4(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G8gat), .B(G36gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n344_), .A2(new_n350_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n344_), .B2(new_n350_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n358_), .A2(KEYINPUT27), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n339_), .A2(new_n342_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n347_), .A2(KEYINPUT20), .A3(new_n349_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(new_n342_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n357_), .B1(new_n355_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT27), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n302_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n272_), .A2(new_n274_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n327_), .A2(new_n328_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(new_n283_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT79), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT31), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n368_), .B(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G71gat), .B(G99gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT30), .ZN(new_n374_));
  XOR2_X1   g173(.A(G15gat), .B(G43gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n372_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n274_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n273_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n344_), .A2(new_n350_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n355_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n291_), .A2(new_n292_), .A3(new_n299_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n299_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n355_), .A2(new_n382_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n362_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT95), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n362_), .A2(new_n390_), .A3(new_n387_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT96), .B1(new_n386_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n384_), .B2(KEYINPUT33), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n291_), .A2(KEYINPUT33), .A3(new_n292_), .A4(new_n299_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n396_), .A2(new_n358_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT94), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n227_), .A2(new_n285_), .ZN(new_n399_));
  AOI211_X1 g198(.A(new_n218_), .B(new_n283_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n288_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n401_), .B2(new_n299_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n284_), .A2(new_n289_), .A3(new_n286_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT94), .A3(new_n297_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n300_), .A2(KEYINPUT93), .A3(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n395_), .A2(new_n397_), .A3(new_n406_), .A4(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n389_), .A2(new_n391_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n301_), .A2(new_n410_), .A3(new_n411_), .A4(new_n383_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n393_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n366_), .B(new_n377_), .C1(new_n380_), .C2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n377_), .A2(new_n301_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n359_), .A2(new_n364_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n415_), .B(new_n416_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT73), .B(G22gat), .ZN(new_n419_));
  INV_X1    g218(.A(G15gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G1gat), .ZN(new_n422_));
  INV_X1    g221(.A(G8gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G1gat), .B(G8gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G29gat), .B(G36gat), .ZN(new_n428_));
  INV_X1    g227(.A(G43gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G50gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n431_), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  NAND2_X1  g235(.A1(G229gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n431_), .B(KEYINPUT15), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n427_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n432_), .A2(KEYINPUT75), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT75), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n437_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n439_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G141gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(new_n320_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(new_n241_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n448_), .B(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n418_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT97), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT98), .ZN(new_n457_));
  AND2_X1   g256(.A1(G230gat), .A2(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT68), .ZN(new_n459_));
  INV_X1    g258(.A(G57gat), .ZN(new_n460_));
  INV_X1    g259(.A(G64gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G57gat), .A2(G64gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G71gat), .A2(G78gat), .ZN(new_n466_));
  INV_X1    g265(.A(G71gat), .ZN(new_n467_));
  INV_X1    g266(.A(G78gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT67), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n462_), .A2(new_n464_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT67), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n465_), .A2(new_n475_), .A3(new_n466_), .A4(new_n469_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n471_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n459_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n473_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(KEYINPUT68), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G85gat), .B(G92gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT9), .ZN(new_n486_));
  AND3_X1   g285(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n486_), .B(new_n489_), .C1(KEYINPUT9), .C2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n492_), .A2(KEYINPUT64), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT64), .B1(new_n492_), .B2(new_n493_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n491_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n501_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT65), .A3(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n500_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n485_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(KEYINPUT66), .A3(new_n485_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(KEYINPUT8), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n500_), .A2(new_n489_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n485_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n496_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n484_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n484_), .A2(new_n517_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n458_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT12), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n484_), .B2(new_n517_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n458_), .B1(new_n484_), .B2(new_n517_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n496_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n508_), .A2(KEYINPUT66), .A3(new_n485_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT66), .B1(new_n508_), .B2(new_n485_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n515_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n516_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n525_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n477_), .A2(new_n478_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT12), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(new_n524_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n521_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(new_n247_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n321_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n521_), .A2(new_n533_), .A3(new_n538_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT69), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT16), .B(G183gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G211gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G127gat), .B(G155gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT68), .B1(new_n554_), .B2(KEYINPUT17), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(new_n427_), .Z(new_n556_));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(new_n531_), .Z(new_n559_));
  NOR2_X1   g358(.A1(new_n554_), .A2(KEYINPUT17), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n431_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n517_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  OAI221_X1 g364(.A(new_n563_), .B1(KEYINPUT35), .B2(new_n565_), .C1(new_n440_), .C2(new_n517_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n441_), .A2(new_n530_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n569_), .A2(KEYINPUT35), .A3(new_n565_), .A4(new_n563_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(G134gat), .ZN(new_n572_));
  INV_X1    g371(.A(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT36), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n568_), .A2(new_n570_), .B1(new_n579_), .B2(new_n574_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT37), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT72), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n568_), .A2(new_n570_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n574_), .A2(new_n579_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n577_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT71), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n584_), .B1(new_n590_), .B2(new_n582_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT71), .B1(new_n587_), .B2(new_n577_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n592_), .A2(KEYINPUT70), .A3(KEYINPUT72), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n583_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT72), .B1(new_n592_), .B2(KEYINPUT70), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n588_), .B2(KEYINPUT70), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n561_), .B1(new_n594_), .B2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n456_), .A2(new_n457_), .A3(new_n550_), .A4(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n454_), .A2(new_n455_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT97), .B1(new_n418_), .B2(new_n453_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n550_), .B(new_n600_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT98), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n601_), .A2(new_n605_), .A3(new_n422_), .A4(new_n301_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n561_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n550_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n453_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n581_), .B(KEYINPUT100), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n418_), .B2(new_n615_), .ZN(new_n616_));
  AOI211_X1 g415(.A(KEYINPUT101), .B(new_n614_), .C1(new_n414_), .C2(new_n417_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n609_), .B(new_n612_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n302_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n606_), .A2(new_n607_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n608_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(G1324gat));
  OAI21_X1  g422(.A(G8gat), .B1(new_n618_), .B2(new_n416_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT103), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(G8gat), .C1(new_n618_), .C2(new_n416_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(KEYINPUT39), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n416_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n601_), .A2(new_n605_), .A3(new_n423_), .A4(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n624_), .A2(KEYINPUT103), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n628_), .A2(new_n635_), .A3(new_n630_), .A4(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(KEYINPUT40), .A3(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n618_), .B2(new_n377_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT41), .Z(new_n643_));
  AND2_X1   g442(.A1(new_n601_), .A2(new_n605_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n377_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n420_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(G1326gat));
  INV_X1    g446(.A(new_n380_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(G22gat), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT106), .Z(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G22gat), .B1(new_n618_), .B2(new_n648_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT105), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT105), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(KEYINPUT42), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT42), .B1(new_n653_), .B2(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  AND2_X1   g456(.A1(new_n456_), .A2(new_n550_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n615_), .A2(new_n609_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n301_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n591_), .A2(new_n593_), .A3(new_n583_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n598_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n418_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n561_), .A3(new_n612_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n671_), .B2(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n302_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n662_), .B1(new_n674_), .B2(G29gat), .ZN(G1328gat));
  OAI21_X1  g474(.A(G36gat), .B1(new_n673_), .B2(new_n416_), .ZN(new_n676_));
  INV_X1    g475(.A(G36gat), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n658_), .A2(new_n677_), .A3(new_n629_), .A4(new_n659_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n678_), .A2(new_n679_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n676_), .A2(KEYINPUT46), .A3(new_n680_), .A4(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1329gat));
  XOR2_X1   g485(.A(KEYINPUT109), .B(G43gat), .Z(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n660_), .B2(new_n377_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n670_), .A2(G43gat), .A3(new_n672_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n377_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g490(.A(G50gat), .B1(new_n661_), .B2(new_n380_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n670_), .A2(G50gat), .A3(new_n672_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n380_), .ZN(G1331gat));
  NOR2_X1   g493(.A1(new_n550_), .A2(new_n453_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n609_), .B(new_n695_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT111), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(G57gat), .A3(new_n301_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n418_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n600_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT110), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n301_), .B1(new_n701_), .B2(KEYINPUT110), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n460_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n698_), .A2(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(new_n701_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n461_), .A3(new_n629_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n697_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G64gat), .B1(new_n708_), .B2(new_n416_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT48), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT48), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1333gat));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n467_), .A3(new_n645_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G71gat), .B1(new_n708_), .B2(new_n377_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(KEYINPUT49), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(KEYINPUT49), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(G1334gat));
  NAND3_X1  g516(.A1(new_n706_), .A2(new_n468_), .A3(new_n380_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G78gat), .B1(new_n708_), .B2(new_n648_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT50), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT50), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(G1335gat));
  NOR3_X1   g521(.A1(new_n699_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n301_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n667_), .A2(new_n561_), .A3(new_n695_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n302_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n726_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n723_), .B2(new_n629_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n725_), .A2(new_n416_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g529(.A(G99gat), .B1(new_n725_), .B2(new_n377_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n723_), .A2(new_n645_), .A3(new_n492_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n723_), .A2(new_n493_), .A3(new_n380_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n667_), .A2(new_n561_), .A3(new_n380_), .A4(new_n695_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(G106gat), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n737_), .B2(G106gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(KEYINPUT112), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n737_), .A2(G106gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n739_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n744_), .B1(new_n747_), .B2(new_n736_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n735_), .B1(new_n743_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n742_), .A2(KEYINPUT112), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n744_), .A3(new_n736_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(KEYINPUT53), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1339gat));
  INV_X1    g552(.A(KEYINPUT119), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n446_), .A2(KEYINPUT117), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n444_), .B(new_n756_), .C1(new_n445_), .C2(new_n442_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n438_), .A3(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n451_), .C1(new_n438_), .C2(new_n436_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n448_), .A2(new_n452_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n542_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n523_), .A2(new_n524_), .A3(new_n532_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n523_), .A2(new_n532_), .A3(new_n518_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n763_), .A2(KEYINPUT55), .B1(new_n458_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n533_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT114), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n533_), .A2(new_n769_), .A3(new_n766_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n765_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT115), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n765_), .A2(new_n768_), .A3(new_n773_), .A4(new_n770_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n539_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n539_), .A4(new_n774_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n775_), .A2(KEYINPUT116), .A3(new_n776_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n453_), .A3(new_n541_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n762_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n615_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(KEYINPUT57), .A3(new_n615_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n777_), .A2(new_n788_), .A3(new_n779_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n775_), .A2(KEYINPUT118), .A3(new_n776_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n541_), .A3(new_n761_), .A4(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n790_), .A2(new_n541_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(KEYINPUT58), .A3(new_n761_), .A4(new_n789_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n795_), .A3(new_n665_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n786_), .A2(new_n787_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n561_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n546_), .A2(new_n453_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n609_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n600_), .A2(new_n804_), .A3(new_n805_), .A4(new_n799_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n754_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT119), .B(new_n807_), .C1(new_n797_), .C2(new_n561_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n416_), .A2(new_n301_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n380_), .A2(new_n377_), .A3(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814_), .B2(new_n453_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(G113gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n798_), .A2(new_n808_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n813_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n811_), .A2(new_n813_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n817_), .B(new_n820_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n822_));
  OAI21_X1  g621(.A(G113gat), .B1(new_n611_), .B2(new_n816_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n815_), .B1(new_n822_), .B2(new_n823_), .ZN(G1340gat));
  OAI21_X1  g623(.A(new_n275_), .B1(new_n550_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n814_), .B(new_n825_), .C1(KEYINPUT60), .C2(new_n275_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n550_), .B(new_n820_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n275_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n814_), .B2(new_n609_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n561_), .B(new_n820_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n814_), .B2(new_n614_), .ZN(new_n832_));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n833_), .B(new_n820_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n834_), .B2(new_n665_), .ZN(G1343gat));
  INV_X1    g634(.A(new_n812_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n648_), .A2(new_n645_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n811_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n838_), .A2(G141gat), .A3(new_n611_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G141gat), .B1(new_n838_), .B2(new_n611_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1344gat));
  OR3_X1    g640(.A1(new_n838_), .A2(G148gat), .A3(new_n550_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G148gat), .B1(new_n838_), .B2(new_n550_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1345gat));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n838_), .A2(new_n561_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n838_), .B2(new_n561_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1346gat));
  INV_X1    g649(.A(new_n665_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n838_), .A2(new_n573_), .A3(new_n851_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n838_), .A2(new_n615_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n573_), .B2(new_n853_), .ZN(G1347gat));
  NOR3_X1   g653(.A1(new_n416_), .A2(new_n301_), .A3(new_n377_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n818_), .A2(new_n648_), .A3(new_n453_), .A4(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n320_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n856_), .B(new_n857_), .C1(KEYINPUT123), .C2(KEYINPUT62), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n856_), .A2(new_n311_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n860_), .A2(new_n862_), .A3(new_n861_), .A4(KEYINPUT124), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1348gat));
  NAND3_X1  g666(.A1(new_n818_), .A2(new_n648_), .A3(new_n855_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n310_), .B1(new_n869_), .B2(new_n610_), .ZN(new_n870_));
  AND4_X1   g669(.A1(G176gat), .A2(new_n811_), .A3(new_n648_), .A4(new_n610_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n855_), .ZN(G1349gat));
  NAND4_X1  g671(.A1(new_n811_), .A2(new_n609_), .A3(new_n648_), .A4(new_n855_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n609_), .A2(new_n331_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n873_), .A2(new_n304_), .B1(new_n869_), .B2(new_n874_), .ZN(G1350gat));
  NOR2_X1   g674(.A1(new_n868_), .A2(new_n851_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n614_), .A2(new_n314_), .ZN(new_n877_));
  OAI22_X1  g676(.A1(new_n876_), .A2(new_n305_), .B1(new_n868_), .B2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT125), .ZN(G1351gat));
  NAND2_X1  g678(.A1(new_n837_), .A2(new_n302_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT126), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n416_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT127), .B1(new_n811_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n884_), .A2(new_n453_), .A3(new_n541_), .A4(new_n781_), .ZN(new_n885_));
  AOI211_X1 g684(.A(new_n785_), .B(new_n614_), .C1(new_n885_), .C2(new_n762_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n783_), .B2(new_n615_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n609_), .B1(new_n888_), .B2(new_n796_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT119), .B1(new_n889_), .B2(new_n807_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n798_), .A2(new_n754_), .A3(new_n808_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(KEYINPUT127), .A4(new_n882_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n453_), .B1(new_n883_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G197gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n891_), .A3(new_n882_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n892_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n241_), .A3(new_n453_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n900_), .ZN(G1352gat));
  AOI21_X1  g700(.A(G204gat), .B1(new_n899_), .B2(new_n610_), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n247_), .B(new_n550_), .C1(new_n898_), .C2(new_n892_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1353gat));
  OR2_X1    g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n899_), .B2(new_n609_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n561_), .B(new_n907_), .C1(new_n898_), .C2(new_n892_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1354gat));
  AOI21_X1  g708(.A(G218gat), .B1(new_n899_), .B2(new_n614_), .ZN(new_n910_));
  INV_X1    g709(.A(G218gat), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n911_), .B(new_n851_), .C1(new_n898_), .C2(new_n892_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1355gat));
endmodule


