//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  INV_X1    g007(.A(G43gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G50gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT15), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT15), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT7), .ZN(new_n221_));
  OAI22_X1  g020(.A1(new_n220_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .A4(KEYINPUT65), .ZN(new_n226_));
  AND4_X1   g025(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  AND2_X1   g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  INV_X1    g031(.A(G92gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G85gat), .A2(G92gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT8), .B1(new_n227_), .B2(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n231_), .A2(new_n236_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .A4(new_n226_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT8), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT9), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n216_), .A2(new_n218_), .B1(new_n229_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G99gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n224_), .A2(KEYINPUT10), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n225_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n234_), .A2(KEYINPUT9), .A3(new_n235_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n245_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT64), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n245_), .A2(new_n249_), .A3(new_n253_), .A4(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n213_), .A2(new_n214_), .B1(new_n243_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n241_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n252_), .A2(new_n254_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n258_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n243_), .A2(KEYINPUT67), .A3(new_n255_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT73), .B1(new_n265_), .B2(new_n212_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267_));
  INV_X1    g066(.A(new_n212_), .ZN(new_n268_));
  AOI211_X1 g067(.A(new_n267_), .B(new_n268_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n207_), .B(new_n257_), .C1(new_n266_), .C2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n204_), .A2(new_n206_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n243_), .A2(KEYINPUT67), .A3(new_n255_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT67), .B1(new_n243_), .B2(new_n255_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n212_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n267_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(KEYINPUT73), .A3(new_n212_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n256_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n271_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n207_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G190gat), .B(G218gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G134gat), .ZN(new_n282_));
  INV_X1    g081(.A(G162gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT75), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n272_), .A2(new_n280_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n284_), .B(KEYINPUT36), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n272_), .B2(new_n280_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT37), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n289_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n270_), .A2(new_n271_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n279_), .B1(new_n278_), .B2(new_n207_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n290_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n292_), .A2(KEYINPUT76), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n289_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n295_), .B1(new_n302_), .B2(KEYINPUT37), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G155gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT16), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G183gat), .ZN(new_n306_));
  INV_X1    g105(.A(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G64gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G71gat), .B(G78gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n313_));
  XOR2_X1   g112(.A(G71gat), .B(G78gat), .Z(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(KEYINPUT11), .A3(new_n309_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G15gat), .B(G22gat), .ZN(new_n319_));
  INV_X1    g118(.A(G1gat), .ZN(new_n320_));
  INV_X1    g119(.A(G8gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT14), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G8gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n318_), .B(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n308_), .B1(new_n327_), .B2(KEYINPUT77), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n328_), .B(KEYINPUT17), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n308_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n303_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT1), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(G155gat), .A3(G162gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n337_), .B(new_n338_), .C1(new_n342_), .C2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n338_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n336_), .B2(KEYINPUT89), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT89), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n353_), .B2(KEYINPUT90), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n336_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n350_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n340_), .A2(new_n341_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n343_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n348_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n362_));
  AND2_X1   g161(.A1(G127gat), .A2(G134gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G127gat), .A2(G134gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G127gat), .ZN(new_n366_));
  INV_X1    g165(.A(G134gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G127gat), .A2(G134gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT87), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G113gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n365_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n373_));
  INV_X1    g172(.A(G120gat), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n363_), .A2(new_n364_), .A3(new_n362_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT87), .B1(new_n368_), .B2(new_n369_), .ZN(new_n377_));
  OAI21_X1  g176(.A(G113gat), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n365_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n379_));
  AOI21_X1  g178(.A(G120gat), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n361_), .B1(new_n375_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n374_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(G120gat), .A3(new_n379_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n352_), .A2(new_n353_), .B1(new_n336_), .B2(new_n356_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n359_), .B(new_n343_), .C1(new_n384_), .C2(new_n350_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .A4(new_n348_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n381_), .A2(new_n386_), .A3(KEYINPUT97), .A4(KEYINPUT4), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n381_), .A2(KEYINPUT4), .A3(new_n386_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT97), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n381_), .B2(KEYINPUT4), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n387_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT0), .ZN(new_n397_));
  INV_X1    g196(.A(G57gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n381_), .A2(new_n386_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n393_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n394_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT33), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n399_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n381_), .A2(new_n393_), .A3(new_n386_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT25), .B(G183gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(G190gat), .ZN(new_n416_));
  INV_X1    g215(.A(G190gat), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n417_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n413_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(KEYINPUT80), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G190gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n415_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n412_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT24), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427_));
  MUX2_X1   g226(.A(new_n426_), .B(KEYINPUT24), .S(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(G183gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT23), .B1(new_n429_), .B2(new_n417_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT23), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(G183gat), .A3(G190gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n421_), .A2(G190gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n417_), .A2(KEYINPUT80), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT26), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT81), .B1(new_n417_), .B2(KEYINPUT26), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n414_), .A2(new_n415_), .A3(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n436_), .A2(KEYINPUT82), .A3(new_n439_), .A4(new_n413_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n424_), .A2(new_n428_), .A3(new_n433_), .A4(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n432_), .A2(KEYINPUT84), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n430_), .A2(new_n432_), .A3(KEYINPUT84), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n429_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G176gat), .ZN(new_n446_));
  AND2_X1   g245(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n449_), .A2(KEYINPUT83), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(KEYINPUT83), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n445_), .A2(new_n450_), .A3(new_n425_), .A4(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G211gat), .B(G218gat), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G197gat), .A2(G204gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT91), .B(G197gat), .ZN(new_n456_));
  OAI211_X1 g255(.A(KEYINPUT21), .B(new_n455_), .C1(new_n456_), .C2(G204gat), .ZN(new_n457_));
  INV_X1    g256(.A(G197gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT92), .B1(new_n458_), .B2(G204gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460_));
  INV_X1    g259(.A(G204gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(G197gat), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n459_), .B(new_n462_), .C1(new_n456_), .C2(new_n461_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n454_), .B(new_n457_), .C1(new_n463_), .C2(KEYINPUT21), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(KEYINPUT21), .A3(new_n453_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n441_), .A2(new_n452_), .A3(new_n464_), .A4(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n433_), .B1(G183gat), .B2(G190gat), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n449_), .A2(KEYINPUT94), .A3(new_n425_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT94), .B1(new_n449_), .B2(new_n425_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT26), .B(G190gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n413_), .A2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n428_), .A2(new_n472_), .A3(new_n443_), .A4(new_n442_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n464_), .A2(new_n465_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n466_), .A2(new_n476_), .A3(KEYINPUT20), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n478_), .B(KEYINPUT93), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT19), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n470_), .A2(new_n464_), .A3(new_n473_), .A4(new_n465_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n441_), .A2(new_n452_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT95), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n441_), .A2(new_n452_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n475_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n484_), .A4(new_n483_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n481_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT96), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G8gat), .B(G36gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT18), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G64gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G92gat), .ZN(new_n497_));
  INV_X1    g296(.A(G64gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n495_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n233_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n492_), .A2(new_n493_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n493_), .B1(new_n492_), .B2(new_n501_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n492_), .A2(new_n501_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n408_), .A2(new_n411_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(new_n500_), .A3(KEYINPUT32), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n481_), .A2(new_n491_), .A3(new_n487_), .A4(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n399_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n382_), .A2(new_n383_), .B1(new_n385_), .B2(new_n348_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT97), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n381_), .A2(KEYINPUT4), .A3(new_n386_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n392_), .B1(new_n516_), .B2(new_n387_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n511_), .B1(new_n517_), .B2(new_n401_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n403_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n507_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(KEYINPUT99), .A2(KEYINPUT20), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT99), .A2(KEYINPUT20), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n484_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT100), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT100), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n484_), .A2(new_n526_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n489_), .A3(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n528_), .A2(new_n480_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n477_), .A2(new_n480_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n520_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n510_), .A2(new_n519_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n506_), .A2(new_n532_), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n361_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT28), .B1(new_n361_), .B2(KEYINPUT29), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G228gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(G22gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n536_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n361_), .A2(KEYINPUT29), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n475_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(G50gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G78gat), .B(G106gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n543_), .A2(new_n544_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n540_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n540_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n543_), .A2(new_n544_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n545_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT101), .B1(new_n533_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT101), .ZN(new_n555_));
  AOI211_X1 g354(.A(new_n555_), .B(new_n552_), .C1(new_n506_), .C2(new_n532_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n382_), .A2(new_n383_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT86), .B(G15gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G71gat), .B(G99gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G227gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT31), .B(G43gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n488_), .B(new_n567_), .Z(new_n568_));
  XOR2_X1   g367(.A(new_n562_), .B(new_n568_), .Z(new_n569_));
  NOR2_X1   g368(.A1(new_n553_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(new_n552_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n505_), .A2(KEYINPUT27), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n501_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n504_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(KEYINPUT27), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n519_), .B(KEYINPUT102), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OAI22_X1  g380(.A1(new_n557_), .A2(new_n569_), .B1(new_n573_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n316_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n265_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n316_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n585_));
  OAI211_X1 g384(.A(G230gat), .B(G233gat), .C1(new_n584_), .C2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT68), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G176gat), .B(G204gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G120gat), .B(G148gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n265_), .B2(new_n583_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n585_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597_));
  OAI211_X1 g396(.A(KEYINPUT12), .B(new_n316_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(new_n586_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n588_), .B(new_n593_), .C1(new_n600_), .C2(new_n587_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n593_), .B(KEYINPUT70), .Z(new_n602_));
  AOI21_X1  g401(.A(new_n587_), .B1(new_n599_), .B2(new_n586_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n586_), .A2(new_n587_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(KEYINPUT71), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(KEYINPUT71), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT79), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n212_), .B(KEYINPUT15), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n326_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n268_), .A2(new_n326_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n212_), .B(new_n325_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n618_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625_));
  INV_X1    g424(.A(G169gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(new_n458_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n621_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n629_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n615_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n630_), .A3(KEYINPUT79), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n614_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n582_), .A2(new_n637_), .ZN(new_n638_));
  NOR4_X1   g437(.A1(new_n335_), .A2(G1gat), .A3(new_n638_), .A4(new_n580_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT104), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(KEYINPUT104), .ZN(new_n643_));
  INV_X1    g442(.A(new_n636_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n606_), .A2(new_n608_), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n601_), .A2(new_n605_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n331_), .B(new_n644_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT103), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n613_), .A2(new_n649_), .A3(new_n331_), .A4(new_n644_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n292_), .A2(KEYINPUT76), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n299_), .B(new_n291_), .C1(new_n272_), .C2(new_n280_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n288_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n651_), .A2(new_n654_), .A3(new_n582_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n580_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .A4(new_n657_), .ZN(G1324gat));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n321_), .B1(new_n655_), .B2(new_n578_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(KEYINPUT106), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(KEYINPUT106), .B2(new_n660_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n333_), .B(KEYINPUT78), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n663_), .A2(new_n321_), .A3(new_n637_), .A4(new_n582_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT105), .B1(new_n664_), .B2(new_n579_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n335_), .A2(new_n638_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n321_), .A4(new_n578_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n660_), .A2(KEYINPUT106), .A3(KEYINPUT39), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n662_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n662_), .A2(new_n669_), .A3(new_n670_), .A4(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  INV_X1    g474(.A(G15gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n666_), .A2(new_n676_), .A3(new_n569_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n655_), .A2(new_n569_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n678_), .B2(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1326gat));
  NAND3_X1  g480(.A1(new_n666_), .A2(new_n538_), .A3(new_n552_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n651_), .A2(new_n582_), .A3(new_n654_), .A4(new_n552_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G22gat), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT107), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(new_n686_), .A3(G22gat), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n685_), .A2(KEYINPUT42), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT42), .B1(new_n685_), .B2(new_n687_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n682_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1327gat));
  NAND2_X1  g491(.A1(new_n302_), .A2(new_n332_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n638_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(G29gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n580_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n637_), .A2(new_n332_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT110), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n303_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n295_), .B(KEYINPUT109), .C1(new_n302_), .C2(KEYINPUT37), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n702_), .B1(new_n706_), .B2(new_n582_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n406_), .B1(new_n405_), .B2(new_n399_), .ZN(new_n708_));
  NOR4_X1   g507(.A1(new_n517_), .A2(KEYINPUT33), .A3(new_n511_), .A4(new_n401_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n492_), .A2(new_n501_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT96), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n492_), .A2(new_n493_), .A3(new_n501_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n576_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n411_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n710_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n532_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n553_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n555_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n533_), .A2(KEYINPUT101), .A3(new_n553_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n573_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n578_), .A2(new_n696_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n721_), .A2(new_n571_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n303_), .A2(new_n702_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n699_), .B(new_n701_), .C1(new_n707_), .C2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n704_), .A2(new_n705_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n728_), .B2(new_n724_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n726_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n698_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n696_), .B(new_n727_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n733_), .A2(KEYINPUT111), .A3(G29gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT111), .B1(new_n733_), .B2(G29gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n697_), .B1(new_n734_), .B2(new_n735_), .ZN(G1328gat));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n578_), .B(new_n727_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(G36gat), .ZN(new_n739_));
  INV_X1    g538(.A(G36gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n693_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n582_), .A2(new_n740_), .A3(new_n637_), .A4(new_n741_), .ZN(new_n742_));
  OR3_X1    g541(.A1(new_n742_), .A2(KEYINPUT112), .A3(new_n579_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT112), .B1(new_n742_), .B2(new_n579_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(KEYINPUT45), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n737_), .B1(new_n739_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n738_), .A2(G36gat), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n751_), .A2(KEYINPUT46), .A3(new_n748_), .A4(new_n747_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1329gat));
  OAI21_X1  g552(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n569_), .A2(G43gat), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n209_), .A2(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n694_), .A2(new_n569_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G43gat), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n754_), .A2(new_n755_), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g560(.A(G50gat), .B1(new_n754_), .B2(new_n553_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n694_), .A2(new_n211_), .A3(new_n552_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n613_), .A2(new_n644_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n582_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n663_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n398_), .B1(new_n767_), .B2(new_n580_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT114), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n654_), .A3(new_n331_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n770_), .A2(new_n398_), .A3(new_n580_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1332gat));
  OAI21_X1  g571(.A(G64gat), .B1(new_n770_), .B2(new_n579_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT48), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n578_), .A2(new_n498_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n767_), .B2(new_n775_), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n770_), .B2(new_n571_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT49), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n571_), .A2(G71gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n767_), .B2(new_n779_), .ZN(G1334gat));
  OAI21_X1  g579(.A(G78gat), .B1(new_n770_), .B2(new_n553_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT50), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n553_), .A2(G78gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n767_), .B2(new_n783_), .ZN(G1335gat));
  OAI211_X1 g583(.A(new_n332_), .B(new_n765_), .C1(new_n707_), .C2(new_n726_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(new_n232_), .A3(new_n580_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n766_), .A2(new_n741_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n766_), .A2(KEYINPUT115), .A3(new_n741_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n696_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n793_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n786_), .B1(new_n794_), .B2(new_n795_), .ZN(G1336gat));
  NOR3_X1   g595(.A1(new_n785_), .A2(new_n233_), .A3(new_n579_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n791_), .A2(new_n578_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n233_), .ZN(G1337gat));
  OAI211_X1 g598(.A(new_n791_), .B(new_n569_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G99gat), .B1(new_n785_), .B2(new_n571_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT51), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n804_), .A3(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1338gat));
  XNOR2_X1  g605(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n807_));
  OAI21_X1  g606(.A(G106gat), .B1(new_n785_), .B2(new_n553_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT52), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(G106gat), .C1(new_n785_), .C2(new_n553_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n552_), .A2(new_n225_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n807_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n807_), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n817_), .B(new_n814_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n617_), .A2(new_n623_), .A3(new_n620_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n622_), .A2(new_n618_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n628_), .A3(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n630_), .A2(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n606_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n595_), .A2(new_n598_), .A3(new_n596_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AND3_X1   g627(.A1(KEYINPUT120), .A2(G230gat), .A3(G233gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n599_), .B2(new_n827_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n826_), .A2(new_n827_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n829_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n602_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n835_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n644_), .A2(new_n601_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n825_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n820_), .B1(new_n840_), .B2(new_n302_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n644_), .A2(new_n601_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n837_), .B2(new_n836_), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT57), .B(new_n654_), .C1(new_n843_), .C2(new_n825_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT122), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n601_), .A2(new_n824_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n601_), .A2(KEYINPUT121), .A3(new_n824_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n838_), .A2(new_n847_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n847_), .B1(new_n838_), .B2(new_n852_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n294_), .B1(new_n654_), .B2(new_n293_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n332_), .B1(new_n845_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n636_), .A2(new_n331_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n859_), .A2(new_n855_), .A3(new_n613_), .A4(new_n860_), .ZN(new_n861_));
  OR2_X1    g660(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n857_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n578_), .A2(new_n580_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n572_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT123), .Z(new_n867_));
  AND2_X1   g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n644_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n864_), .A2(new_n870_), .A3(new_n867_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n636_), .A2(new_n371_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n869_), .B1(new_n873_), .B2(new_n874_), .ZN(G1340gat));
  OAI21_X1  g674(.A(new_n374_), .B1(new_n613_), .B2(KEYINPUT60), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n868_), .B(new_n876_), .C1(KEYINPUT60), .C2(new_n374_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n871_), .A2(new_n872_), .A3(new_n613_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n374_), .ZN(G1341gat));
  AOI21_X1  g678(.A(G127gat), .B1(new_n868_), .B2(new_n331_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n332_), .A2(new_n366_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n873_), .B2(new_n881_), .ZN(G1342gat));
  AOI21_X1  g681(.A(G134gat), .B1(new_n868_), .B2(new_n302_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n855_), .A2(new_n367_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n873_), .B2(new_n884_), .ZN(G1343gat));
  INV_X1    g684(.A(new_n570_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n857_), .B2(new_n863_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(new_n865_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n644_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n614_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n331_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n888_), .B2(new_n302_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n728_), .A2(new_n283_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n888_), .B2(new_n897_), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n579_), .A2(new_n696_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n569_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n553_), .ZN(new_n903_));
  AOI211_X1 g702(.A(new_n901_), .B(new_n903_), .C1(new_n857_), .C2(new_n863_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n626_), .B1(new_n904_), .B2(new_n644_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n905_), .A2(KEYINPUT62), .ZN(new_n906_));
  INV_X1    g705(.A(new_n901_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n903_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n864_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n447_), .A2(new_n448_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n909_), .A2(new_n636_), .A3(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT62), .B1(new_n911_), .B2(new_n905_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n906_), .A2(new_n912_), .ZN(G1348gat));
  NAND2_X1  g712(.A1(new_n904_), .A2(new_n614_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g714(.A1(new_n909_), .A2(new_n332_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n413_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n429_), .B2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n909_), .B2(new_n855_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n904_), .A2(new_n302_), .A3(new_n471_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1351gat));
  INV_X1    g720(.A(new_n899_), .ZN(new_n922_));
  AOI211_X1 g721(.A(new_n886_), .B(new_n922_), .C1(new_n857_), .C2(new_n863_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n644_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n887_), .A2(new_n899_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n613_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(KEYINPUT125), .B2(new_n461_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT125), .B(G204gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1353gat));
  AOI21_X1  g729(.A(new_n332_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n931_), .A2(KEYINPUT126), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(KEYINPUT126), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n923_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  OR2_X1    g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1354gat));
  INV_X1    g735(.A(G218gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n926_), .B2(new_n654_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n303_), .A2(G218gat), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n938_), .B(new_n939_), .C1(new_n926_), .C2(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G218gat), .B1(new_n923_), .B2(new_n302_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n926_), .A2(new_n940_), .ZN(new_n943_));
  OAI21_X1  g742(.A(KEYINPUT127), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n941_), .A2(new_n944_), .ZN(G1355gat));
endmodule


