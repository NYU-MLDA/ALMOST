//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT81), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n203_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT31), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G227gat), .A2(G233gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT80), .Z(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT78), .B(G169gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT79), .ZN(new_n218_));
  OR2_X1    g017(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n219_));
  INV_X1    g018(.A(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(new_n223_), .A3(KEYINPUT23), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n213_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(G183gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n220_), .A2(KEYINPUT26), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G190gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(KEYINPUT77), .B(new_n230_), .C1(new_n234_), .C2(new_n239_), .ZN(new_n240_));
  NOR3_X1   g039(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n219_), .A2(KEYINPUT25), .A3(new_n221_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT26), .B(G190gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n235_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT77), .B1(new_n246_), .B2(new_n230_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n226_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT30), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G15gat), .B(G43gat), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n226_), .B(KEYINPUT30), .C1(new_n243_), .C2(new_n247_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n250_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n210_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G71gat), .B(G99gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n253_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n230_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT30), .B1(new_n262_), .B2(new_n226_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n251_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n210_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n250_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n256_), .A2(new_n257_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n257_), .B1(new_n256_), .B2(new_n267_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n208_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n256_), .A2(new_n267_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n257_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n275_), .A2(new_n269_), .A3(new_n268_), .A4(new_n207_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(KEYINPUT83), .A3(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OR3_X1    g080(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283_));
  INV_X1    g082(.A(G141gat), .ZN(new_n284_));
  INV_X1    g083(.A(G148gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n282_), .A2(new_n286_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n290_));
  INV_X1    g089(.A(G155gat), .ZN(new_n291_));
  INV_X1    g090(.A(G162gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n289_), .A2(new_n293_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(KEYINPUT1), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G155gat), .A3(G162gat), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n293_), .A2(new_n297_), .A3(new_n299_), .A4(new_n294_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G141gat), .B(G148gat), .Z(new_n301_));
  AND3_X1   g100(.A1(new_n300_), .A2(KEYINPUT85), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT85), .B1(new_n300_), .B2(new_n301_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n296_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT86), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n306_), .B(new_n296_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(G197gat), .A2(G204gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G197gat), .A2(G204gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT87), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT21), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n314_), .ZN(new_n316_));
  INV_X1    g115(.A(G218gat), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n317_), .A2(G211gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(G211gat), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n318_), .A2(new_n319_), .B1(new_n312_), .B2(new_n311_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n315_), .B1(new_n321_), .B2(KEYINPUT21), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G228gat), .A2(G233gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(KEYINPUT21), .ZN(new_n325_));
  INV_X1    g124(.A(new_n315_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(KEYINPUT29), .B2(new_n304_), .ZN(new_n328_));
  OAI22_X1  g127(.A1(new_n310_), .A2(new_n324_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G78gat), .B(G106gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G22gat), .B(G50gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n308_), .A2(new_n334_), .A3(new_n309_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(new_n335_), .A3(new_n332_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n331_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n340_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT88), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n331_), .A3(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n203_), .B(new_n204_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n305_), .A2(new_n350_), .A3(new_n307_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n302_), .A2(new_n303_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n206_), .A2(new_n352_), .A3(new_n296_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT4), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n351_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n354_), .A2(new_n356_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n360_), .B2(new_n367_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n349_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n360_), .A2(new_n367_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n365_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(KEYINPUT95), .A3(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n327_), .B1(new_n262_), .B2(new_n226_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT19), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n241_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n385_));
  INV_X1    g184(.A(G183gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT25), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .A4(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n385_), .A2(new_n218_), .A3(new_n224_), .A4(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT22), .B(G169gat), .ZN(new_n390_));
  INV_X1    g189(.A(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n215_), .A2(new_n217_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n229_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT20), .B1(new_n322_), .B2(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n382_), .A2(new_n384_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n384_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n262_), .A2(new_n327_), .A3(new_n226_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n322_), .B2(new_n396_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n381_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n402_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n384_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n381_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n389_), .A2(new_n395_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n401_), .B1(new_n327_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n248_), .A2(new_n322_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n399_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n404_), .A2(KEYINPUT90), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT27), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n411_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT90), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n381_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT97), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT97), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n413_), .A2(new_n417_), .A3(new_n420_), .A4(new_n414_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n412_), .A2(KEYINPUT27), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n384_), .B1(new_n382_), .B2(new_n397_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n400_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n407_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n422_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n428_), .A2(KEYINPUT96), .A3(KEYINPUT27), .A4(new_n412_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n419_), .A2(new_n421_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n348_), .A2(new_n376_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n413_), .A2(new_n417_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n357_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n366_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n434_));
  OR2_X1    g233(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n435_));
  OAI221_X1 g234(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .C1(new_n370_), .C2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n370_), .A2(new_n435_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n407_), .A2(KEYINPUT32), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT94), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n439_), .B(new_n443_), .ZN(new_n444_));
  OAI22_X1  g243(.A1(new_n444_), .A2(new_n415_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n445_));
  AOI211_X1 g244(.A(new_n442_), .B(new_n445_), .C1(new_n373_), .C2(new_n368_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n347_), .B1(new_n438_), .B2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n281_), .B1(new_n431_), .B2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n272_), .A2(new_n276_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(new_n375_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT98), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n430_), .A2(new_n451_), .ZN(new_n452_));
  AOI221_X4 g251(.A(KEYINPUT98), .B1(new_n427_), .B2(new_n429_), .C1(new_n419_), .C2(new_n421_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n450_), .B(new_n347_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT99), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n419_), .A2(new_n421_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n427_), .A2(new_n429_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT98), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n430_), .A2(new_n451_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(KEYINPUT99), .A3(new_n347_), .A4(new_n450_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n448_), .B1(new_n456_), .B2(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G29gat), .B(G36gat), .Z(new_n465_));
  XOR2_X1   g264(.A(G43gat), .B(G50gat), .Z(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(KEYINPUT15), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT74), .B(G8gat), .ZN(new_n470_));
  INV_X1    g269(.A(G1gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G8gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n469_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n476_), .A2(new_n467_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT75), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n476_), .B(new_n467_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n480_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n479_), .A2(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G113gat), .B(G141gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(G169gat), .B(G197gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n464_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n495_));
  XOR2_X1   g294(.A(G71gat), .B(G78gat), .Z(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n495_), .A2(new_n496_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(new_n476_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504_));
  XOR2_X1   g303(.A(G127gat), .B(G155gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT16), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G183gat), .B(G211gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(KEYINPUT17), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n513_));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT6), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  OR3_X1    g319(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G85gat), .B(G92gat), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT67), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n524_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT10), .B(G99gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT64), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT65), .B(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT66), .B(G92gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT9), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(G85gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n523_), .A2(KEYINPUT9), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n532_), .A2(new_n535_), .A3(new_n536_), .A4(new_n519_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n528_), .A2(new_n537_), .ZN(new_n538_));
  OAI221_X1 g337(.A(new_n516_), .B1(KEYINPUT71), .B2(new_n517_), .C1(new_n538_), .C2(new_n467_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT68), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n528_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n537_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n542_), .B2(new_n469_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n517_), .A2(KEYINPUT71), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G134gat), .B(G162gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT36), .Z(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n543_), .B(new_n544_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT37), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(KEYINPUT73), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n551_), .A2(new_n553_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n545_), .A2(new_n561_), .A3(new_n549_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .A4(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n512_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n542_), .A2(KEYINPUT12), .A3(new_n499_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n499_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n528_), .B2(new_n537_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT12), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n538_), .A2(new_n499_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n565_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(G230gat), .B(G233gat), .C1(new_n570_), .C2(new_n568_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G120gat), .B(G148gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT69), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n577_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n580_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT13), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT13), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n580_), .B1(new_n581_), .B2(new_n577_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n582_), .B1(KEYINPUT69), .B2(new_n579_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n564_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n492_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n471_), .A3(new_n375_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n589_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n595_), .A2(new_n491_), .A3(new_n512_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n456_), .A2(new_n463_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n448_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n558_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n376_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n592_), .A2(new_n593_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n602_), .A3(new_n603_), .ZN(G1324gat));
  INV_X1    g403(.A(new_n462_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n591_), .A2(new_n605_), .A3(new_n470_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT100), .Z(new_n607_));
  OAI21_X1  g406(.A(G8gat), .B1(new_n601_), .B2(new_n462_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT39), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g410(.A(new_n281_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G15gat), .B1(new_n601_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT101), .Z(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(KEYINPUT41), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(KEYINPUT41), .ZN(new_n616_));
  INV_X1    g415(.A(new_n591_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n617_), .A2(G15gat), .A3(new_n612_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n601_), .B2(new_n347_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n347_), .A2(G22gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n617_), .B2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n512_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n600_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n589_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n492_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n628_), .A2(G29gat), .A3(new_n376_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n595_), .A2(new_n491_), .A3(new_n624_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n557_), .A2(new_n563_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT43), .B1(new_n464_), .B2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n464_), .A2(KEYINPUT43), .A3(new_n631_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  INV_X1    g435(.A(new_n631_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n599_), .A2(new_n634_), .A3(new_n636_), .A4(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n630_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT103), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n640_), .A2(KEYINPUT103), .A3(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT44), .B(new_n630_), .C1(new_n635_), .C2(new_n639_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(new_n375_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(KEYINPUT104), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G29gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT104), .B1(new_n645_), .B2(new_n647_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n629_), .B1(new_n649_), .B2(new_n650_), .ZN(G1328gat));
  XNOR2_X1  g450(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n646_), .A2(new_n605_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n599_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT102), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n638_), .A3(new_n632_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n654_), .B(KEYINPUT44), .C1(new_n657_), .C2(new_n630_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n653_), .B1(new_n658_), .B2(new_n642_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  INV_X1    g459(.A(G36gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n627_), .A2(new_n661_), .A3(new_n605_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n652_), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n652_), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n664_), .B(new_n667_), .C1(new_n659_), .C2(G36gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1329gat));
  INV_X1    g468(.A(G43gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n449_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n646_), .B(new_n671_), .C1(new_n658_), .C2(new_n642_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n628_), .B2(new_n612_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT47), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n676_), .A3(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n627_), .B2(new_n348_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n645_), .A2(new_n646_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n348_), .A2(G50gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(G1331gat));
  NOR2_X1   g481(.A1(new_n512_), .A2(new_n490_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n599_), .A2(new_n595_), .A3(new_n600_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(G57gat), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n376_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n599_), .A2(KEYINPUT106), .A3(new_n491_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(new_n464_), .B2(new_n490_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n687_), .A2(new_n595_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n564_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n376_), .B1(new_n691_), .B2(KEYINPUT107), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(KEYINPUT107), .B2(new_n691_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n686_), .B1(new_n693_), .B2(new_n685_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n684_), .B2(new_n462_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT108), .Z(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT48), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(KEYINPUT48), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n691_), .A2(G64gat), .A3(new_n462_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(G1333gat));
  OR3_X1    g499(.A1(new_n691_), .A2(G71gat), .A3(new_n612_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G71gat), .B1(new_n684_), .B2(new_n612_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT109), .ZN(G1334gat));
  OAI21_X1  g504(.A(G78gat), .B1(new_n684_), .B2(new_n347_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT50), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n347_), .A2(G78gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT110), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n691_), .B2(new_n709_), .ZN(G1335gat));
  INV_X1    g509(.A(G85gat), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n589_), .A2(new_n490_), .A3(new_n624_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n657_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT111), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n657_), .A2(new_n715_), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n711_), .B1(new_n717_), .B2(new_n375_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n690_), .A2(new_n625_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n719_), .A2(G85gat), .A3(new_n376_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1336gat));
  NAND3_X1  g520(.A1(new_n717_), .A2(new_n605_), .A3(new_n533_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n719_), .A2(new_n462_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(G92gat), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT112), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n722_), .B(new_n726_), .C1(G92gat), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1337gat));
  NAND4_X1  g527(.A1(new_n690_), .A2(new_n277_), .A3(new_n530_), .A4(new_n625_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n612_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n730_));
  INV_X1    g529(.A(G99gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n657_), .A2(new_n348_), .A3(new_n712_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G106gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G106gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n348_), .A2(new_n531_), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n736_), .A2(new_n737_), .B1(new_n719_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g539(.A1(new_n490_), .A2(new_n579_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n565_), .A2(new_n571_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT55), .B1(new_n744_), .B2(new_n566_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n572_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n744_), .A2(KEYINPUT55), .A3(new_n566_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT56), .B1(new_n748_), .B2(new_n577_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n750_), .B(new_n578_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n743_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n477_), .A2(new_n478_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n481_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n754_), .B2(new_n753_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n487_), .B1(new_n482_), .B2(new_n481_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n756_), .A2(new_n757_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n583_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n752_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n600_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(KEYINPUT117), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n764_));
  INV_X1    g563(.A(new_n600_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n752_), .B2(new_n759_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(KEYINPUT57), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(KEYINPUT57), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n579_), .A2(new_n758_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT58), .B(new_n769_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n637_), .A3(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n763_), .A2(new_n767_), .A3(new_n768_), .A4(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n564_), .A2(new_n491_), .A3(new_n589_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n564_), .A2(new_n491_), .A3(new_n589_), .A4(new_n777_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(KEYINPUT114), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(KEYINPUT114), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n512_), .A2(new_n775_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n348_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n376_), .A2(new_n449_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT118), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n775_), .A2(new_n512_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n782_), .A2(new_n783_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  INV_X1    g591(.A(new_n787_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n788_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(G113gat), .B1(new_n795_), .B2(new_n490_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n768_), .A2(new_n774_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n766_), .A2(KEYINPUT57), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n512_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT59), .B(new_n787_), .C1(new_n790_), .C2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(KEYINPUT59), .C1(new_n784_), .C2(new_n787_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n800_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n490_), .A2(G113gat), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT120), .Z(new_n808_));
  AOI21_X1  g607(.A(new_n796_), .B1(new_n806_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n589_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n795_), .B(new_n811_), .C1(KEYINPUT60), .C2(new_n810_), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n589_), .B(new_n800_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n810_), .ZN(G1341gat));
  XNOR2_X1  g613(.A(KEYINPUT122), .B(G127gat), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n624_), .A2(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n816_), .B(new_n800_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n788_), .A2(new_n794_), .A3(new_n624_), .ZN(new_n818_));
  INV_X1    g617(.A(G127gat), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT121), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n817_), .B1(new_n821_), .B2(new_n823_), .ZN(G1342gat));
  AOI21_X1  g623(.A(G134gat), .B1(new_n795_), .B2(new_n765_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT123), .B(G134gat), .Z(new_n826_));
  NOR2_X1   g625(.A1(new_n631_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n806_), .B2(new_n827_), .ZN(G1343gat));
  NAND4_X1  g627(.A1(new_n462_), .A2(new_n612_), .A3(new_n348_), .A4(new_n375_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT124), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n791_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n491_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(new_n284_), .ZN(G1344gat));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n589_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n285_), .ZN(G1345gat));
  NOR2_X1   g634(.A1(new_n831_), .A2(new_n512_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT61), .B(G155gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  OAI21_X1  g637(.A(G162gat), .B1(new_n831_), .B2(new_n631_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n765_), .A2(new_n292_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n831_), .B2(new_n840_), .ZN(G1347gat));
  AOI21_X1  g640(.A(new_n348_), .B1(new_n790_), .B2(new_n799_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n462_), .A2(new_n612_), .A3(new_n375_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n490_), .A3(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n845_));
  INV_X1    g644(.A(new_n390_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n844_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT62), .B1(new_n844_), .B2(G169gat), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1348gat));
  NAND2_X1  g648(.A1(new_n842_), .A2(new_n843_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n391_), .B1(new_n850_), .B2(new_n589_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n784_), .A2(new_n348_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(G176gat), .A3(new_n595_), .A4(new_n843_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1349gat));
  AND2_X1   g653(.A1(new_n235_), .A2(new_n387_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n843_), .A2(new_n624_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n842_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n852_), .A2(new_n857_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT125), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n231_), .A2(new_n232_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(G1350gat));
  OAI21_X1  g661(.A(G190gat), .B1(new_n850_), .B2(new_n631_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n765_), .A2(new_n245_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n850_), .B2(new_n864_), .ZN(G1351gat));
  INV_X1    g664(.A(KEYINPUT126), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n462_), .A2(new_n281_), .A3(new_n347_), .A4(new_n375_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n791_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n490_), .ZN(new_n870_));
  INV_X1    g669(.A(G197gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n866_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n871_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n869_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n490_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(G1352gat));
  NOR2_X1   g674(.A1(new_n868_), .A2(new_n589_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT127), .B(G204gat), .Z(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n876_), .B2(new_n879_), .ZN(G1353gat));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n868_), .A2(new_n512_), .A3(new_n881_), .A4(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n869_), .A2(new_n624_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n881_), .ZN(G1354gat));
  OAI21_X1  g684(.A(G218gat), .B1(new_n868_), .B2(new_n631_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n765_), .A2(new_n317_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n868_), .B2(new_n887_), .ZN(G1355gat));
endmodule


