//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_,
    new_n972_, new_n973_, new_n974_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n998_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT92), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT31), .B(G15gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G71gat), .B(G99gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G43gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n205_), .B(new_n207_), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT85), .B(G183gat), .Z(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT25), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT85), .B(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT25), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT86), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT87), .B(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(G183gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n212_), .A2(new_n215_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n227_), .A2(KEYINPUT88), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(G176gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n235_), .A2(new_n229_), .A3(new_n228_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT88), .B1(new_n227_), .B2(new_n231_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n222_), .A2(new_n232_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT30), .ZN(new_n240_));
  INV_X1    g039(.A(new_n235_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT22), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT89), .B1(new_n242_), .B2(G169gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G169gat), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n234_), .B(new_n243_), .C1(new_n244_), .C2(KEYINPUT89), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n210_), .A2(new_n219_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n224_), .A2(KEYINPUT90), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT90), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n241_), .B(new_n245_), .C1(new_n246_), .C2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n239_), .A2(new_n240_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n240_), .B1(new_n239_), .B2(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT91), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n252_), .A2(KEYINPUT91), .A3(new_n253_), .ZN(new_n256_));
  INV_X1    g055(.A(G127gat), .ZN(new_n257_));
  INV_X1    g056(.A(G134gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G127gat), .A2(G134gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G113gat), .ZN(new_n262_));
  INV_X1    g061(.A(G113gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n262_), .A2(G120gat), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(G120gat), .B1(new_n262_), .B2(new_n264_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n255_), .A2(new_n256_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n252_), .A2(KEYINPUT91), .A3(new_n253_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(new_n254_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n209_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n267_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n254_), .A3(new_n269_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n208_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n272_), .A2(new_n275_), .A3(KEYINPUT93), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT93), .B1(new_n272_), .B2(new_n275_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G78gat), .B(G106gat), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G228gat), .A2(G233gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT97), .Z(new_n282_));
  NOR2_X1   g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT1), .Z(new_n288_));
  OR2_X1    g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G141gat), .ZN(new_n292_));
  INV_X1    g091(.A(G148gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT94), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT3), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n283_), .A2(KEYINPUT94), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n285_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n295_), .A2(new_n297_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n289_), .A2(new_n287_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n301_), .A2(KEYINPUT95), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT95), .B1(new_n301_), .B2(new_n302_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n291_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n306_));
  XOR2_X1   g105(.A(G197gat), .B(G204gat), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT21), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n307_), .B2(KEYINPUT21), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n309_), .B(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n282_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n281_), .A2(KEYINPUT97), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n311_), .B(new_n308_), .ZN(new_n315_));
  AOI211_X1 g114(.A(new_n314_), .B(new_n315_), .C1(new_n305_), .C2(KEYINPUT29), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n280_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n301_), .A2(new_n302_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n301_), .A2(KEYINPUT95), .A3(new_n302_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n290_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n312_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n282_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n314_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n306_), .A2(new_n312_), .A3(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n279_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G22gat), .B(G50gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT28), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n305_), .A2(KEYINPUT29), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n317_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT98), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n317_), .A2(new_n337_), .A3(new_n329_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT96), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n332_), .B1(new_n305_), .B2(KEYINPUT29), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n322_), .A2(new_n323_), .A3(new_n331_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT96), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n326_), .A2(KEYINPUT98), .A3(new_n279_), .A4(new_n328_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n338_), .A2(new_n346_), .A3(KEYINPUT99), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT99), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n344_), .A2(new_n345_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n317_), .A2(new_n329_), .A3(new_n337_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n336_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT100), .Z(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT19), .Z(new_n356_));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n244_), .A2(new_n234_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n241_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT102), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT102), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n361_), .A3(new_n241_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G183gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n227_), .B1(new_n364_), .B2(new_n217_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n236_), .A2(new_n231_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT25), .B(G183gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT26), .B(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT101), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n369_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n372_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT101), .B1(new_n376_), .B2(new_n368_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n367_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n357_), .B1(new_n378_), .B2(new_n312_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n239_), .A2(new_n250_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n312_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n356_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n312_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n367_), .B(new_n315_), .C1(new_n375_), .C2(new_n377_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT20), .A4(new_n356_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G64gat), .ZN(new_n390_));
  INV_X1    g189(.A(G92gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n383_), .A2(new_n387_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n356_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n365_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n374_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n376_), .A2(KEYINPUT101), .A3(new_n368_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT20), .B1(new_n399_), .B2(new_n315_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n395_), .B1(new_n400_), .B2(new_n381_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n392_), .B1(new_n401_), .B2(new_n386_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n353_), .B1(new_n394_), .B2(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n400_), .A2(new_n395_), .A3(new_n381_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n369_), .A2(new_n373_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n312_), .A2(new_n396_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n315_), .B1(new_n239_), .B2(new_n250_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n356_), .B1(new_n408_), .B2(KEYINPUT20), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n393_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n401_), .A2(new_n392_), .A3(new_n386_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(KEYINPUT27), .A3(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n403_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n305_), .A2(new_n269_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n267_), .B(new_n291_), .C1(new_n304_), .C2(new_n303_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(KEYINPUT4), .A3(new_n415_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n305_), .A2(new_n269_), .A3(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G85gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT0), .ZN(new_n426_));
  INV_X1    g225(.A(G57gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n418_), .B2(new_n423_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n352_), .A2(new_n413_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n401_), .A2(new_n386_), .A3(new_n434_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n436_), .B(new_n437_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n429_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n393_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n418_), .A2(new_n423_), .A3(KEYINPUT33), .A4(new_n428_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n411_), .A4(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n419_), .A2(new_n417_), .A3(new_n422_), .ZN(new_n444_));
  AOI211_X1 g243(.A(new_n428_), .B(new_n444_), .C1(new_n420_), .C2(new_n416_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n438_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n336_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT99), .B1(new_n338_), .B2(new_n346_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n349_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n278_), .B1(new_n433_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n272_), .A2(new_n275_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n403_), .A2(new_n412_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n432_), .ZN(new_n456_));
  NOR4_X1   g255(.A1(new_n352_), .A2(new_n454_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G120gat), .B(G148gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT5), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(G176gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(G204gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(G204gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(KEYINPUT67), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n462_), .A2(KEYINPUT67), .A3(new_n463_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G230gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G85gat), .B(G92gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT9), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(G99gat), .A3(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(G99gat), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n479_), .A2(KEYINPUT10), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(KEYINPUT10), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n478_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n391_), .A2(KEYINPUT9), .ZN(new_n483_));
  OR2_X1    g282(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n472_), .A2(new_n477_), .A3(new_n482_), .A4(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI211_X1 g290(.A(KEYINPUT8), .B(new_n470_), .C1(new_n491_), .C2(new_n477_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(new_n479_), .A3(new_n478_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n475_), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n488_), .B(new_n495_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n493_), .B1(new_n498_), .B2(new_n471_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n487_), .B1(new_n492_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT11), .ZN(new_n501_));
  INV_X1    g300(.A(G64gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n427_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G57gat), .A2(G64gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  INV_X1    g307(.A(G71gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G78gat), .ZN(new_n510_));
  INV_X1    g309(.A(G78gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G71gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n507_), .A2(new_n508_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n508_), .B1(new_n507_), .B2(new_n513_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n506_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n504_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G57gat), .A2(G64gat), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT11), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G71gat), .B(G78gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT65), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n507_), .A2(new_n508_), .A3(new_n513_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n505_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n469_), .B1(new_n500_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n500_), .A2(new_n524_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n500_), .A2(new_n524_), .A3(KEYINPUT12), .ZN(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT66), .B(new_n469_), .C1(new_n500_), .C2(new_n524_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(new_n530_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n500_), .A2(new_n524_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n528_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n469_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n468_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n538_), .A2(new_n465_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT13), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n543_), .B(new_n544_), .C1(new_n468_), .C2(new_n539_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT84), .ZN(new_n548_));
  XOR2_X1   g347(.A(G169gat), .B(G197gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(G50gat), .ZN(new_n554_));
  INV_X1    g353(.A(G29gat), .ZN(new_n555_));
  INV_X1    g354(.A(G36gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT68), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G29gat), .A2(G36gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n558_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n561_), .A2(G43gat), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(G43gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G29gat), .B(G36gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT68), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n566_), .B2(new_n560_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n554_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G43gat), .B1(new_n561_), .B2(new_n562_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n564_), .A3(new_n560_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(G50gat), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  INV_X1    g372(.A(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G8gat), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n572_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT15), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n572_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n568_), .A2(KEYINPUT15), .A3(new_n571_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n582_), .B1(new_n586_), .B2(new_n581_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n582_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n572_), .A2(new_n581_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n548_), .B(new_n553_), .C1(new_n589_), .C2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n553_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n592_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(KEYINPUT84), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n458_), .A2(new_n547_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT81), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n603_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT80), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT75), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n579_), .A2(new_n580_), .A3(new_n612_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n523_), .A3(new_n516_), .A4(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n524_), .B1(new_n617_), .B2(new_n613_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n608_), .A2(new_n609_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n609_), .B1(new_n608_), .B2(new_n619_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(KEYINPUT76), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT76), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n616_), .A2(new_n618_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n623_), .A2(new_n606_), .A3(new_n625_), .A4(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n599_), .B1(new_n622_), .B2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n627_), .B(KEYINPUT81), .C1(new_n620_), .C2(new_n621_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n598_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(G134gat), .ZN(new_n634_));
  INV_X1    g433(.A(G162gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT36), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT71), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT34), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT35), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n572_), .A2(new_n500_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n500_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT69), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n585_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT15), .B1(new_n568_), .B2(new_n571_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n500_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT69), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n641_), .B1(new_n646_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n640_), .B(KEYINPUT35), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n644_), .A2(new_n642_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n638_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n641_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n642_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n656_), .B1(new_n649_), .B2(KEYINPUT69), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n644_), .A2(new_n645_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n653_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT36), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n636_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT70), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n660_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n654_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT74), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT74), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n654_), .A2(new_n664_), .A3(new_n668_), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n586_), .A2(new_n645_), .A3(new_n500_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n650_), .A2(new_n671_), .A3(new_n656_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n653_), .B1(new_n672_), .B2(new_n655_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n638_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT72), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT72), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n638_), .C1(new_n651_), .C2(new_n653_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n664_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT37), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n670_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n632_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n574_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT38), .ZN(new_n684_));
  OAI22_X1  g483(.A1(new_n683_), .A2(new_n432_), .B1(KEYINPUT105), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(KEYINPUT38), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n622_), .A2(new_n628_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n654_), .A2(new_n664_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT103), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n654_), .A2(new_n664_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n598_), .A2(new_n688_), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT104), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G1gat), .B1(new_n697_), .B2(new_n432_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT105), .B(new_n684_), .C1(new_n683_), .C2(new_n432_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n687_), .A2(new_n698_), .A3(new_n699_), .ZN(G1324gat));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n695_), .A2(new_n413_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n575_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT106), .B(G8gat), .C1(new_n695_), .C2(new_n413_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(KEYINPUT39), .A3(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n682_), .A2(new_n575_), .A3(new_n455_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT39), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n701_), .B(new_n707_), .C1(new_n702_), .C2(new_n575_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1325gat));
  INV_X1    g510(.A(new_n682_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n278_), .ZN(new_n713_));
  OR3_X1    g512(.A1(new_n712_), .A2(G15gat), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G15gat), .B1(new_n697_), .B2(new_n713_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n716_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1326gat));
  OR3_X1    g518(.A1(new_n712_), .A2(G22gat), .A3(new_n450_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G22gat), .B1(new_n697_), .B2(new_n450_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT42), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT42), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(G1327gat));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(KEYINPUT44), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n681_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(KEYINPUT43), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(KEYINPUT43), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n681_), .B(new_n731_), .C1(new_n452_), .C2(new_n457_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n729_), .A2(new_n730_), .A3(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n593_), .A2(new_n596_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n631_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n546_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT107), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n726_), .B1(new_n734_), .B2(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n450_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n446_), .A2(new_n450_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n713_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n457_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n680_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT108), .B1(new_n744_), .B2(new_n731_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n727_), .A2(new_n728_), .A3(KEYINPUT43), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n732_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n726_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n738_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n739_), .A2(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n751_), .A2(new_n555_), .A3(new_n432_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n694_), .A2(new_n631_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n598_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G29gat), .B1(new_n755_), .B2(new_n456_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n752_), .A2(new_n756_), .ZN(G1328gat));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n556_), .A3(new_n455_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT45), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n748_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n413_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(new_n556_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n759_), .B(KEYINPUT46), .C1(new_n762_), .C2(new_n556_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1329gat));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n454_), .A2(new_n564_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n739_), .A2(new_n750_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771_));
  AOI21_X1  g570(.A(G43gat), .B1(new_n755_), .B2(new_n278_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n770_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n768_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n769_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n760_), .A2(new_n761_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT110), .B1(new_n778_), .B2(new_n772_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n770_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(KEYINPUT47), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n776_), .A2(new_n781_), .ZN(G1330gat));
  OAI21_X1  g581(.A(G50gat), .B1(new_n751_), .B2(new_n450_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n352_), .A2(new_n554_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT111), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n754_), .B2(new_n785_), .ZN(G1331gat));
  NOR3_X1   g585(.A1(new_n458_), .A2(new_n546_), .A3(new_n735_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n631_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n694_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT112), .B1(new_n456_), .B2(G57gat), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n790_), .A2(KEYINPUT112), .A3(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(new_n791_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n788_), .A2(new_n681_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n456_), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n792_), .A2(new_n427_), .B1(new_n793_), .B2(new_n795_), .ZN(G1332gat));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n502_), .A3(new_n455_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n789_), .A2(new_n455_), .A3(new_n694_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT48), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G64gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G64gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT113), .ZN(G1333gat));
  OAI21_X1  g602(.A(G71gat), .B1(new_n790_), .B2(new_n713_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT49), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n794_), .A2(new_n509_), .A3(new_n278_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1334gat));
  NAND3_X1  g606(.A1(new_n794_), .A2(new_n511_), .A3(new_n352_), .ZN(new_n808_));
  OAI21_X1  g607(.A(G78gat), .B1(new_n790_), .B2(new_n450_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT114), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(G78gat), .C1(new_n790_), .C2(new_n450_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n810_), .A2(KEYINPUT50), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT50), .B1(new_n810_), .B2(new_n812_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n808_), .B1(new_n813_), .B2(new_n814_), .ZN(G1335gat));
  NAND2_X1  g614(.A1(new_n787_), .A2(new_n753_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G85gat), .B1(new_n817_), .B2(new_n456_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n546_), .A2(new_n735_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n747_), .A2(new_n736_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n456_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(G1336gat));
  AOI21_X1  g622(.A(G92gat), .B1(new_n817_), .B2(new_n455_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n413_), .A2(new_n391_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n821_), .B2(new_n825_), .ZN(G1337gat));
  OAI21_X1  g625(.A(G99gat), .B1(new_n820_), .B2(new_n713_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n453_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n816_), .B2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g629(.A1(new_n817_), .A2(new_n478_), .A3(new_n352_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n747_), .A2(new_n352_), .A3(new_n736_), .A4(new_n819_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G106gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G106gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g636(.A1(new_n352_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n456_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n688_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n842_));
  AND3_X1   g641(.A1(new_n533_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n533_), .B2(new_n842_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n500_), .A2(new_n524_), .A3(KEYINPUT12), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT12), .B1(new_n500_), .B2(new_n524_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n847_), .A2(KEYINPUT55), .A3(new_n527_), .A4(new_n532_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n530_), .A2(new_n534_), .A3(new_n531_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n536_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n843_), .A2(new_n844_), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n468_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  INV_X1    g653(.A(new_n468_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n533_), .A2(new_n842_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT118), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n533_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n854_), .B(new_n855_), .C1(new_n859_), .C2(new_n851_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n853_), .A2(new_n543_), .A3(new_n735_), .A4(new_n860_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n587_), .A2(new_n588_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n590_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n553_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n595_), .B2(new_n553_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n694_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT120), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n693_), .B1(new_n861_), .B2(new_n866_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(KEYINPUT57), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n868_), .A2(new_n875_), .A3(new_n869_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT119), .B1(new_n871_), .B2(KEYINPUT57), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n853_), .A2(new_n865_), .A3(new_n543_), .A4(new_n860_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT58), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n681_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n840_), .B1(new_n879_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n631_), .A2(new_n597_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n885_), .A2(new_n886_), .B1(new_n545_), .B2(new_n542_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n631_), .A2(KEYINPUT115), .A3(new_n597_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n680_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT116), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n680_), .A2(new_n887_), .A3(new_n891_), .A4(new_n888_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n890_), .A2(KEYINPUT54), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT54), .B1(new_n890_), .B2(new_n892_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n839_), .B1(new_n884_), .B2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G113gat), .B1(new_n896_), .B2(new_n735_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n868_), .A2(new_n869_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n873_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n872_), .B1(new_n871_), .B2(KEYINPUT57), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n882_), .B(new_n900_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n736_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n899_), .B1(new_n895_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n839_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n870_), .A2(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n688_), .B1(new_n907_), .B2(new_n882_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n894_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n890_), .A2(KEYINPUT54), .A3(new_n892_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n906_), .B1(new_n908_), .B2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n905_), .B1(new_n912_), .B2(KEYINPUT59), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n597_), .A2(new_n263_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n897_), .B1(new_n913_), .B2(new_n914_), .ZN(G1340gat));
  XNOR2_X1  g714(.A(KEYINPUT121), .B(G120gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n913_), .B2(new_n547_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n546_), .B2(KEYINPUT60), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n917_), .A2(KEYINPUT60), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n896_), .A2(new_n919_), .A3(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT122), .B1(new_n918_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n905_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n924_), .B(new_n547_), .C1(new_n896_), .C2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n916_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n928_), .A3(new_n921_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n923_), .A2(new_n929_), .ZN(G1341gat));
  AOI21_X1  g729(.A(G127gat), .B1(new_n896_), .B2(new_n631_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n840_), .A2(new_n257_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n913_), .B2(new_n932_), .ZN(G1342gat));
  OAI21_X1  g732(.A(new_n258_), .B1(new_n912_), .B2(new_n694_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n924_), .B1(new_n896_), .B2(new_n925_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n680_), .A2(new_n258_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n934_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(KEYINPUT123), .B(new_n934_), .C1(new_n935_), .C2(new_n937_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1343gat));
  NOR2_X1   g741(.A1(new_n450_), .A2(new_n455_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n278_), .A2(new_n432_), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n943_), .B(new_n944_), .C1(new_n908_), .C2(new_n911_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n597_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n292_), .ZN(G1344gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n546_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n293_), .ZN(G1345gat));
  NOR2_X1   g748(.A1(new_n945_), .A2(new_n736_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT61), .B(G155gat), .Z(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1346gat));
  NOR3_X1   g751(.A1(new_n945_), .A2(new_n635_), .A3(new_n680_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n635_), .B1(new_n945_), .B2(new_n694_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n954_), .A2(KEYINPUT124), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(KEYINPUT124), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n953_), .B1(new_n955_), .B2(new_n956_), .ZN(G1347gat));
  NOR2_X1   g756(.A1(new_n413_), .A2(new_n456_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n713_), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  AOI211_X1 g760(.A(new_n352_), .B(new_n961_), .C1(new_n895_), .C2(new_n904_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n233_), .B1(new_n962_), .B2(new_n735_), .ZN(new_n963_));
  OR2_X1    g762(.A1(new_n963_), .A2(KEYINPUT62), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n962_), .A2(new_n735_), .A3(new_n244_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(KEYINPUT62), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n964_), .A2(new_n965_), .A3(new_n966_), .ZN(G1348gat));
  AOI21_X1  g766(.A(G176gat), .B1(new_n962_), .B2(new_n547_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n908_), .A2(new_n911_), .ZN(new_n969_));
  NOR4_X1   g768(.A1(new_n969_), .A2(new_n234_), .A3(new_n546_), .A4(new_n352_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n968_), .B1(new_n960_), .B2(new_n970_), .ZN(G1349gat));
  INV_X1    g770(.A(new_n962_), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n972_), .A2(new_n840_), .A3(new_n370_), .ZN(new_n973_));
  OR4_X1    g772(.A1(new_n352_), .A2(new_n969_), .A3(new_n736_), .A4(new_n961_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n974_), .B2(new_n210_), .ZN(G1350gat));
  OAI21_X1  g774(.A(G190gat), .B1(new_n972_), .B2(new_n680_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n962_), .A2(new_n371_), .A3(new_n693_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1351gat));
  NOR2_X1   g777(.A1(new_n278_), .A2(new_n450_), .ZN(new_n979_));
  OAI211_X1 g778(.A(new_n958_), .B(new_n979_), .C1(new_n908_), .C2(new_n911_), .ZN(new_n980_));
  INV_X1    g779(.A(new_n980_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n981_), .A2(new_n735_), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n982_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g782(.A1(new_n980_), .A2(new_n546_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  XOR2_X1   g785(.A(KEYINPUT125), .B(G204gat), .Z(new_n987_));
  OAI21_X1  g786(.A(new_n986_), .B1(new_n984_), .B2(new_n987_), .ZN(G1353gat));
  OAI22_X1  g787(.A1(new_n980_), .A2(new_n840_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n989_));
  AOI21_X1  g788(.A(new_n959_), .B1(new_n884_), .B2(new_n895_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(KEYINPUT63), .B(G211gat), .ZN(new_n991_));
  NAND4_X1  g790(.A1(new_n990_), .A2(new_n688_), .A3(new_n979_), .A4(new_n991_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n989_), .A2(new_n992_), .ZN(new_n993_));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994_));
  XNOR2_X1  g793(.A(new_n993_), .B(new_n994_), .ZN(G1354gat));
  XNOR2_X1  g794(.A(KEYINPUT127), .B(G218gat), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n980_), .A2(new_n680_), .A3(new_n996_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n981_), .A2(new_n693_), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n997_), .B1(new_n998_), .B2(new_n996_), .ZN(G1355gat));
endmodule


