//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .A4(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G57gat), .B(G64gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT11), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G71gat), .B(G78gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n214_), .A2(KEYINPUT11), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(KEYINPUT11), .B2(new_n214_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n218_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n209_), .A2(KEYINPUT65), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n208_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT7), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n224_), .B1(new_n232_), .B2(new_n203_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT64), .B(KEYINPUT8), .Z(new_n234_));
  AOI211_X1 g033(.A(new_n202_), .B(new_n234_), .C1(new_n231_), .C2(new_n209_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n213_), .B(new_n223_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n231_), .B1(new_n209_), .B2(KEYINPUT65), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n227_), .A2(new_n228_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n203_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n235_), .B1(new_n241_), .B2(KEYINPUT8), .ZN(new_n242_));
  INV_X1    g041(.A(new_n213_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n222_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(G230gat), .A2(G233gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n222_), .B(KEYINPUT67), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n213_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT12), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n236_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(new_n246_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n244_), .A2(KEYINPUT68), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT68), .B1(new_n244_), .B2(new_n253_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n250_), .B(new_n252_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n247_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G120gat), .B(G148gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT5), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n247_), .A2(new_n256_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT13), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(KEYINPUT13), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT69), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT71), .B(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT72), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n277_), .A3(new_n274_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G1gat), .B(G8gat), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(new_n223_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT73), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n285_), .B(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G127gat), .B(G155gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(G183gat), .B(G211gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n288_), .B1(KEYINPUT17), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT67), .A3(KEYINPUT17), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT37), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G29gat), .B(G36gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT15), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n249_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G232gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT34), .ZN(new_n306_));
  INV_X1    g105(.A(new_n302_), .ZN(new_n307_));
  OAI221_X1 g106(.A(new_n304_), .B1(KEYINPUT35), .B2(new_n306_), .C1(new_n307_), .C2(new_n249_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(KEYINPUT35), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n304_), .B2(KEYINPUT70), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n308_), .B(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G190gat), .B(G218gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT36), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n314_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(KEYINPUT36), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n311_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n299_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n316_), .B(KEYINPUT37), .C1(new_n320_), .C2(new_n311_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n298_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n270_), .A2(KEYINPUT75), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G169gat), .ZN(new_n328_));
  INV_X1    g127(.A(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(KEYINPUT24), .A3(new_n331_), .ZN(new_n332_));
  OR3_X1    g131(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335_));
  INV_X1    g134(.A(G190gat), .ZN(new_n336_));
  OR3_X1    g135(.A1(new_n335_), .A2(new_n336_), .A3(KEYINPUT26), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT25), .B(G183gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT26), .B1(new_n335_), .B2(new_n336_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT23), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n334_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G197gat), .B(G204gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT21), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n349_));
  NOR2_X1   g148(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n350_));
  AND2_X1   g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G197gat), .A2(G204gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n349_), .B(new_n350_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n345_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n348_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n349_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n350_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(KEYINPUT89), .A3(new_n353_), .A4(new_n345_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n347_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n328_), .A2(KEYINPUT22), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G169gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n362_), .B1(new_n364_), .B2(G169gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n329_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n369_), .A2(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT81), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(G176gat), .B1(new_n363_), .B2(new_n362_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G169gat), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n374_), .B(KEYINPUT80), .C1(new_n362_), .C2(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n372_), .A2(new_n376_), .A3(KEYINPUT81), .A4(new_n331_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n342_), .B1(G183gat), .B2(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n343_), .B(new_n361_), .C1(new_n373_), .C2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n356_), .A2(new_n360_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n347_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n338_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT26), .B(G190gat), .Z(new_n386_));
  OAI211_X1 g185(.A(new_n334_), .B(new_n342_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n375_), .A2(KEYINPUT91), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n375_), .A2(KEYINPUT91), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n389_), .A2(new_n390_), .A3(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n378_), .A2(new_n331_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n387_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n381_), .B1(new_n384_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n380_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n378_), .A2(new_n331_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n390_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n388_), .A3(new_n329_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n385_), .A2(new_n386_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n342_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n399_), .A2(new_n401_), .B1(new_n404_), .B2(new_n334_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n381_), .B1(new_n405_), .B2(new_n361_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n397_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n343_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n377_), .A2(new_n378_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n372_), .A2(new_n376_), .A3(new_n331_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n406_), .B(new_n407_), .C1(new_n413_), .C2(new_n361_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT18), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n398_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n395_), .A2(new_n407_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n406_), .B(new_n397_), .C1(new_n413_), .C2(new_n361_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n420_), .A2(new_n423_), .A3(KEYINPUT27), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n412_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n361_), .B1(new_n425_), .B2(new_n343_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n384_), .B2(new_n393_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n426_), .A2(new_n397_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n407_), .B1(new_n380_), .B2(new_n394_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n418_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT27), .B1(new_n430_), .B2(new_n420_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT98), .B1(new_n424_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n428_), .A2(new_n429_), .A3(new_n418_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n419_), .B1(new_n398_), .B2(new_n414_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n420_), .A2(new_n423_), .A3(KEYINPUT27), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n432_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G134gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G127gat), .ZN(new_n442_));
  INV_X1    g241(.A(G127gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G134gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT82), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n444_), .A3(KEYINPUT82), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G113gat), .B(G120gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n447_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n448_), .B1(new_n451_), .B2(new_n445_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G141gat), .A2(G148gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT3), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G141gat), .A2(G148gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT2), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464_));
  AND2_X1   g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(G155gat), .A2(G162gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G155gat), .A2(G162gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT85), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n469_), .A2(KEYINPUT1), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(KEYINPUT1), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G141gat), .B(G148gat), .Z(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n453_), .A2(new_n454_), .A3(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n470_), .A2(new_n467_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n479_), .A2(new_n463_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n481_), .A3(KEYINPUT4), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n453_), .A2(new_n454_), .A3(new_n477_), .A4(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n453_), .A2(new_n477_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n481_), .A2(new_n488_), .A3(new_n483_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT0), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G57gat), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n491_), .A2(KEYINPUT0), .ZN(new_n494_));
  INV_X1    g293(.A(G57gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(KEYINPUT0), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n493_), .A2(new_n497_), .A3(G85gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(G85gat), .B1(new_n493_), .B2(new_n497_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT97), .ZN(new_n502_));
  INV_X1    g301(.A(new_n500_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n487_), .A2(new_n503_), .A3(new_n489_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n502_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT28), .B1(new_n477_), .B2(KEYINPUT29), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT29), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n480_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G22gat), .B(G50gat), .Z(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n513_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G228gat), .A2(G233gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT86), .Z(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT87), .B1(new_n480_), .B2(new_n510_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n361_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n477_), .B2(KEYINPUT29), .ZN(new_n523_));
  INV_X1    g322(.A(new_n519_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n384_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n525_), .A3(KEYINPUT90), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT90), .B1(new_n521_), .B2(new_n525_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G78gat), .B(G106gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  AOI211_X1 g329(.A(KEYINPUT90), .B(new_n530_), .C1(new_n521_), .C2(new_n525_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n517_), .B(new_n526_), .C1(new_n529_), .C2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n521_), .A2(new_n525_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n533_), .B2(KEYINPUT90), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n528_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n517_), .A2(new_n526_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G71gat), .B(G99gat), .ZN(new_n539_));
  INV_X1    g338(.A(G43gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542_));
  INV_X1    g341(.A(G15gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n541_), .B(new_n544_), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT30), .B(new_n343_), .C1(new_n373_), .C2(new_n379_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT30), .B1(new_n425_), .B2(new_n343_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n343_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n453_), .B(KEYINPUT31), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT84), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n555_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n548_), .A2(new_n549_), .A3(new_n546_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n545_), .B1(new_n553_), .B2(new_n547_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT83), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT83), .B(new_n559_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n538_), .B1(new_n558_), .B2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n440_), .A2(new_n507_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n558_), .A2(new_n566_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n504_), .A2(KEYINPUT94), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n481_), .A2(new_n488_), .A3(new_n484_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n500_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n500_), .A2(KEYINPUT95), .A3(new_n575_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n482_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n573_), .B1(new_n504_), .B2(KEYINPUT94), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n430_), .A2(KEYINPUT92), .A3(new_n420_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT92), .B1(new_n430_), .B2(new_n420_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n501_), .A2(new_n504_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n421_), .A2(new_n422_), .A3(KEYINPUT32), .A4(new_n419_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n398_), .A2(new_n414_), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n591_), .A2(KEYINPUT96), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(KEYINPUT96), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n588_), .B(new_n589_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n538_), .B1(new_n587_), .B2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n532_), .B(new_n537_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n596_), .A2(new_n431_), .A3(new_n424_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n572_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n440_), .A2(new_n567_), .A3(KEYINPUT99), .A4(new_n507_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n570_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n269_), .B2(new_n325_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G169gat), .B(G197gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n302_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n276_), .A2(new_n278_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n279_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n307_), .A3(new_n281_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n609_), .A2(KEYINPUT76), .A3(new_n612_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n608_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n608_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n284_), .A2(new_n303_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(new_n609_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n607_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n616_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT76), .B1(new_n609_), .B2(new_n612_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n620_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n606_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT77), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n621_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n621_), .B2(new_n626_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR4_X1   g430(.A1(new_n327_), .A2(new_n601_), .A3(new_n603_), .A4(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n507_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n271_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT38), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n317_), .A2(new_n321_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n268_), .A2(new_n630_), .A3(new_n297_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT101), .A3(new_n600_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT101), .B1(new_n641_), .B2(new_n600_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n507_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n635_), .A2(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n440_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n647_), .A3(new_n600_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n632_), .A2(new_n272_), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n644_), .B2(new_n572_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT41), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(KEYINPUT41), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n632_), .A2(new_n543_), .A3(new_n571_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n632_), .A2(new_n659_), .A3(new_n538_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661_));
  INV_X1    g460(.A(new_n644_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n538_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n663_), .B2(G22gat), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT42), .B(new_n659_), .C1(new_n662_), .C2(new_n538_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n660_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n636_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n297_), .ZN(new_n670_));
  AND4_X1   g469(.A1(new_n600_), .A2(new_n630_), .A3(new_n268_), .A4(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n633_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  INV_X1    g472(.A(new_n268_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(new_n631_), .A3(new_n297_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n600_), .A2(new_n676_), .A3(new_n324_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n600_), .B2(new_n324_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT103), .B(new_n675_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n673_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT104), .B(KEYINPUT44), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n679_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT44), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(G29gat), .A3(new_n633_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n672_), .B1(new_n687_), .B2(new_n690_), .ZN(G1328gat));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n671_), .A2(new_n692_), .A3(new_n647_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT45), .Z(new_n694_));
  OAI211_X1 g493(.A(new_n647_), .B(new_n689_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G36gat), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT105), .B(KEYINPUT46), .Z(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1329gat));
  NAND4_X1  g497(.A1(new_n687_), .A2(G43gat), .A3(new_n571_), .A4(new_n689_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n671_), .A2(new_n571_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n540_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n671_), .A2(new_n704_), .A3(new_n538_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n538_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n688_), .B2(KEYINPUT44), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(KEYINPUT106), .A3(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT106), .B1(new_n708_), .B2(G50gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT107), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n705_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1331gat));
  NOR3_X1   g514(.A1(new_n269_), .A2(new_n601_), .A3(new_n630_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n297_), .A3(new_n669_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n507_), .ZN(new_n718_));
  NOR4_X1   g517(.A1(new_n601_), .A2(new_n326_), .A3(new_n630_), .A4(new_n268_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n495_), .A3(new_n633_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1332gat));
  OAI21_X1  g520(.A(G64gat), .B1(new_n717_), .B2(new_n440_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT48), .ZN(new_n723_));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n724_), .A3(new_n647_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n717_), .B2(new_n572_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  INV_X1    g527(.A(G71gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n719_), .A2(new_n729_), .A3(new_n571_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n717_), .B2(new_n706_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  INV_X1    g532(.A(G78gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n719_), .A2(new_n734_), .A3(new_n538_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1335gat));
  AND2_X1   g535(.A1(new_n716_), .A2(new_n670_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n210_), .A3(new_n633_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n677_), .A2(new_n678_), .ZN(new_n739_));
  NOR4_X1   g538(.A1(new_n739_), .A2(new_n630_), .A3(new_n268_), .A4(new_n297_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n633_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n742_), .B2(new_n210_), .ZN(G1336gat));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n211_), .A3(new_n647_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n740_), .A2(new_n647_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n746_), .B2(new_n211_), .ZN(G1337gat));
  NAND2_X1  g546(.A1(new_n740_), .A2(new_n571_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n571_), .A2(new_n205_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n748_), .A2(G99gat), .B1(new_n737_), .B2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT51), .Z(G1338gat));
  NAND2_X1  g550(.A1(new_n740_), .A2(new_n538_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n206_), .B1(new_n753_), .B2(KEYINPUT109), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(KEYINPUT52), .A3(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n737_), .A2(new_n206_), .A3(new_n538_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT108), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(new_n754_), .B2(new_n756_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT53), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n761_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n757_), .A4(new_n759_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1339gat));
  INV_X1    g565(.A(new_n567_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n647_), .A2(new_n767_), .A3(new_n507_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n256_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n256_), .A2(KEYINPUT112), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n250_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n238_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n246_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n255_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n244_), .A2(KEYINPUT68), .A3(new_n253_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n781_), .A2(KEYINPUT55), .A3(new_n250_), .A4(new_n252_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n778_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n263_), .B1(new_n775_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n769_), .B1(new_n784_), .B2(KEYINPUT113), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(new_n782_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n786_), .B(KEYINPUT56), .C1(new_n788_), .C2(new_n263_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n264_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT111), .B(new_n264_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n785_), .A2(new_n789_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n615_), .A2(new_n608_), .A3(new_n616_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n606_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n619_), .A2(new_n609_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n619_), .A2(KEYINPUT114), .A3(new_n609_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n608_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n796_), .A2(new_n801_), .A3(KEYINPUT115), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n265_), .A2(new_n621_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n636_), .B1(new_n794_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT57), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(KEYINPUT57), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n263_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n784_), .A2(new_n769_), .ZN(new_n812_));
  AND4_X1   g611(.A1(new_n621_), .A2(new_n803_), .A3(new_n264_), .A4(new_n802_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n810_), .B(new_n324_), .C1(new_n814_), .C2(KEYINPUT58), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n324_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n810_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n824_));
  OAI22_X1  g623(.A1(new_n820_), .A2(new_n823_), .B1(new_n805_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT119), .B1(new_n809_), .B2(new_n825_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n822_), .A2(new_n810_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n818_), .B1(new_n822_), .B2(new_n810_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n805_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n824_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n827_), .A2(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n794_), .A2(new_n804_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT57), .A3(new_n669_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT118), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n831_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n297_), .B1(new_n826_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n325_), .A2(new_n631_), .A3(new_n268_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n768_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n630_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n298_), .B1(new_n809_), .B2(new_n825_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n647_), .A2(new_n767_), .A3(KEYINPUT59), .A4(new_n507_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n843_), .A2(KEYINPUT59), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n630_), .A2(G113gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT120), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n845_), .B1(new_n850_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n674_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n844_), .A2(new_n857_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n850_), .A2(new_n270_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n855_), .ZN(G1341gat));
  NAND3_X1  g659(.A1(new_n844_), .A2(new_n443_), .A3(new_n297_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n850_), .A2(new_n297_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n443_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n844_), .B2(new_n636_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n324_), .A2(G134gat), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT121), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n850_), .B2(new_n866_), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n571_), .A2(new_n706_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n869_), .A2(new_n647_), .A3(new_n507_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n831_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n837_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n298_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n874_), .B2(new_n847_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n630_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n270_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n297_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n669_), .A2(G162gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n875_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n875_), .B2(new_n324_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n883_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n839_), .A2(new_n842_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n890_), .A2(new_n821_), .A3(new_n871_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT122), .B(new_n885_), .C1(new_n891_), .C2(new_n887_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(G1347gat));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n440_), .A2(new_n633_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n767_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n848_), .A2(new_n630_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n898_), .B2(G169gat), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n894_), .A3(G169gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n400_), .A2(new_n388_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n901_), .A2(new_n903_), .B1(new_n904_), .B2(new_n898_), .ZN(G1348gat));
  NAND2_X1  g704(.A1(new_n848_), .A2(new_n897_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n329_), .B1(new_n906_), .B2(new_n268_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n896_), .A2(new_n329_), .A3(new_n572_), .A4(new_n538_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n270_), .A2(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n907_), .B1(new_n890_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1349gat));
  NOR2_X1   g711(.A1(new_n906_), .A2(new_n298_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(G183gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n385_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n906_), .B2(new_n821_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n669_), .A2(new_n386_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n906_), .B2(new_n917_), .ZN(G1351gat));
  NOR2_X1   g717(.A1(new_n896_), .A2(new_n869_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n630_), .B(new_n919_), .C1(new_n839_), .C2(new_n842_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT126), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n919_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n874_), .B2(new_n847_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n924_), .A2(KEYINPUT125), .A3(new_n925_), .A4(new_n630_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n922_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(G197gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT125), .B1(new_n924_), .B2(new_n630_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n922_), .B(new_n926_), .C1(new_n931_), .C2(new_n928_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1352gat));
  INV_X1    g732(.A(G204gat), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n924_), .B(new_n270_), .C1(KEYINPUT127), .C2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(KEYINPUT127), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1353gat));
  INV_X1    g736(.A(new_n924_), .ZN(new_n938_));
  OAI22_X1  g737(.A1(new_n938_), .A2(new_n298_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT63), .B(G211gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n924_), .A2(new_n297_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n938_), .B2(new_n821_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n669_), .A2(G218gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n938_), .B2(new_n944_), .ZN(G1355gat));
endmodule


