//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_;
  INV_X1    g000(.A(G204gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT88), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G204gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT87), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n210_), .A3(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT89), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT89), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n206_), .A2(new_n211_), .A3(new_n215_), .A4(new_n212_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G211gat), .B(G218gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT88), .B(G204gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT87), .B(G197gat), .ZN(new_n221_));
  OAI22_X1  g020(.A1(G197gat), .A2(new_n220_), .B1(new_n221_), .B2(G204gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n219_), .B1(new_n222_), .B2(KEYINPUT21), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n218_), .A2(KEYINPUT90), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n206_), .A2(new_n211_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n212_), .B1(new_n218_), .B2(KEYINPUT90), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G228gat), .A2(G233gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n230_), .B(KEYINPUT85), .Z(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT86), .Z(new_n232_));
  XOR2_X1   g031(.A(G155gat), .B(G162gat), .Z(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT83), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236_));
  INV_X1    g035(.A(G141gat), .ZN(new_n237_));
  INV_X1    g036(.A(G148gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .A4(KEYINPUT82), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240_));
  OAI22_X1  g039(.A1(new_n240_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G141gat), .A2(G148gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT2), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n233_), .B1(new_n235_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n233_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n237_), .A2(new_n238_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n242_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n246_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n252_), .A2(KEYINPUT84), .A3(KEYINPUT29), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT84), .B1(new_n252_), .B2(KEYINPUT29), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n229_), .B(new_n232_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n229_), .A2(KEYINPUT92), .ZN(new_n256_));
  INV_X1    g055(.A(new_n228_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT92), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n261_));
  AOI22_X1  g060(.A1(new_n256_), .A2(new_n260_), .B1(new_n252_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n255_), .B1(new_n262_), .B2(new_n231_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n252_), .A2(KEYINPUT29), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT28), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n252_), .A2(new_n261_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n229_), .A2(KEYINPUT92), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n258_), .A2(new_n259_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n231_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n265_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n255_), .A3(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G78gat), .B(G106gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G22gat), .B(G50gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n266_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n266_), .B2(new_n274_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G190gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT26), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT26), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G183gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT25), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G183gat), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n283_), .A2(KEYINPUT79), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n288_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(KEYINPUT24), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT23), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G183gat), .A3(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  OR3_X1    g104(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n300_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n303_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n308_), .B(new_n309_), .C1(G183gat), .C2(G190gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G169gat), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n295_), .A2(new_n307_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G15gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT30), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n313_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n318_), .A2(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT81), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n319_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n325_), .A2(KEYINPUT80), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(KEYINPUT80), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n322_), .B(new_n324_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n317_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G71gat), .B(G99gat), .ZN(new_n330_));
  INV_X1    g129(.A(G43gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT31), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n329_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT100), .ZN(new_n336_));
  XOR2_X1   g135(.A(G1gat), .B(G29gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n322_), .A2(new_n324_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n325_), .B(KEYINPUT80), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT98), .B(KEYINPUT4), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n342_), .A2(new_n252_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT97), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n251_), .B1(new_n233_), .B2(new_n247_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n234_), .B(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n351_), .A2(new_n239_), .A3(new_n244_), .A4(new_n241_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n349_), .B1(new_n352_), .B2(new_n233_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT95), .B1(new_n328_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT95), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n342_), .A2(new_n252_), .A3(new_n355_), .A4(new_n343_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n320_), .A2(new_n325_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT96), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n354_), .A2(new_n356_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n348_), .B1(new_n360_), .B2(KEYINPUT4), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n356_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n353_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n347_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n341_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n364_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n362_), .A2(KEYINPUT4), .A3(new_n363_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n367_), .B(new_n340_), .C1(new_n368_), .C2(new_n348_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n334_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT19), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(G204gat), .B1(new_n208_), .B2(new_n210_), .ZN(new_n378_));
  AOI21_X1  g177(.A(G197gat), .B1(new_n203_), .B2(new_n205_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT21), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n218_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n283_), .A2(new_n285_), .A3(new_n290_), .A4(new_n292_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n383_), .A2(new_n300_), .A3(new_n306_), .A4(new_n305_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n312_), .A2(new_n310_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n228_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n377_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n313_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n373_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n313_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n382_), .B2(new_n257_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n377_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n228_), .A2(new_n385_), .A3(new_n384_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n224_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n395_), .A3(KEYINPUT93), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n224_), .A2(new_n228_), .A3(new_n313_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT20), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n258_), .A2(new_n386_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n375_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n397_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n403_), .B1(new_n397_), .B2(new_n407_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n372_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT102), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n388_), .A2(new_n389_), .A3(new_n373_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT93), .B1(new_n392_), .B2(new_n395_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n407_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n402_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n404_), .B(KEYINPUT20), .C1(new_n258_), .C2(new_n386_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n390_), .A2(new_n396_), .B1(new_n417_), .B2(new_n375_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n403_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(KEYINPUT102), .A3(new_n372_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n412_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT103), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n372_), .B1(new_n418_), .B2(new_n403_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n375_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n256_), .A2(new_n260_), .A3(new_n386_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n389_), .A2(new_n376_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n417_), .A2(new_n375_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n402_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT101), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT101), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n424_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n422_), .A2(new_n423_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n423_), .B1(new_n422_), .B2(new_n435_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n281_), .B(new_n371_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT32), .B(new_n403_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT32), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n418_), .B1(new_n440_), .B2(new_n402_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n370_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n369_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n361_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(KEYINPUT33), .A3(new_n367_), .A4(new_n340_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n340_), .B1(new_n347_), .B2(new_n360_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n345_), .A2(new_n364_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n368_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n442_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n281_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT102), .B1(new_n420_), .B2(new_n372_), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n411_), .B(KEYINPUT27), .C1(new_n416_), .C2(new_n419_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n434_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n433_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n457_));
  OAI22_X1  g256(.A1(new_n454_), .A2(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n266_), .A2(new_n274_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n277_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n278_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n370_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n453_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n334_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n438_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G113gat), .B(G141gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT77), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G169gat), .B(G197gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT15), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT71), .B(KEYINPUT14), .C1(new_n477_), .C2(new_n478_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G8gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n476_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT74), .ZN(new_n488_));
  INV_X1    g287(.A(new_n486_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n487_), .A2(new_n488_), .B1(new_n489_), .B2(new_n475_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n476_), .A2(KEYINPUT74), .A3(new_n486_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT75), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n486_), .B(new_n475_), .Z(new_n495_));
  INV_X1    g294(.A(new_n491_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n490_), .A2(new_n494_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n498_), .A2(KEYINPUT76), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT76), .B1(new_n498_), .B2(new_n499_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n472_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT78), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n471_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n506_), .B(new_n472_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n503_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G120gat), .B(G148gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT5), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G176gat), .B(G204gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(G57gat), .B(G64gat), .Z(new_n516_));
  INV_X1    g315(.A(KEYINPUT11), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n518_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT65), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n525_), .B(KEYINPUT6), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT65), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n528_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G85gat), .B(G92gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n524_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  AOI211_X1 g339(.A(KEYINPUT8), .B(new_n538_), .C1(new_n536_), .C2(new_n529_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT10), .B(G99gat), .Z(new_n543_));
  AOI22_X1  g342(.A1(new_n539_), .A2(KEYINPUT9), .B1(new_n543_), .B2(new_n533_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n544_), .B(new_n529_), .C1(KEYINPUT9), .C2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n523_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n521_), .B(new_n522_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(KEYINPUT12), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n523_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n514_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n513_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n512_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT68), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n553_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n558_), .B2(new_n513_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n512_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n557_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NOR4_X1   g360(.A1(new_n554_), .A2(KEYINPUT68), .A3(new_n555_), .A4(new_n512_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n556_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(KEYINPUT13), .B(new_n556_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n549_), .B(new_n489_), .ZN(new_n569_));
  AND2_X1   g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n571_), .A2(new_n572_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT72), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT73), .B1(new_n571_), .B2(new_n572_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n571_), .A2(KEYINPUT73), .A3(new_n572_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n576_), .B(KEYINPUT17), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n581_), .B(new_n582_), .C1(new_n583_), .C2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT36), .Z(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n542_), .A2(new_n475_), .A3(new_n546_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT69), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  AOI211_X1 g396(.A(KEYINPUT70), .B(new_n597_), .C1(new_n547_), .C2(new_n476_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT35), .A3(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n592_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n590_), .A2(KEYINPUT36), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n605_), .A3(new_n602_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n600_), .A2(new_n605_), .A3(new_n602_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n609_), .B2(new_n603_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n587_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  AND4_X1   g410(.A1(new_n467_), .A2(new_n508_), .A3(new_n568_), .A4(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n477_), .A3(new_n370_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n565_), .A2(new_n508_), .A3(new_n566_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n587_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n565_), .A2(KEYINPUT104), .A3(new_n508_), .A4(new_n566_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n458_), .A2(KEYINPUT103), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n422_), .A2(new_n435_), .A3(new_n423_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n462_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  AOI22_X1  g423(.A1(new_n624_), .A2(new_n371_), .B1(new_n465_), .B2(new_n334_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n609_), .A2(new_n603_), .A3(KEYINPUT105), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT105), .B1(new_n609_), .B2(new_n603_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n621_), .A2(new_n629_), .A3(new_n370_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G1gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n613_), .A2(new_n614_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n615_), .A2(new_n631_), .A3(new_n632_), .ZN(G1324gat));
  NOR2_X1   g432(.A1(new_n436_), .A2(new_n437_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n612_), .A2(new_n478_), .A3(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n621_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(G8gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(G8gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  INV_X1    g441(.A(new_n334_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n612_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n621_), .A2(new_n629_), .A3(new_n643_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(new_n645_), .B2(G15gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT106), .Z(G1326gat));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n612_), .A2(new_n650_), .A3(new_n462_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n621_), .A2(new_n629_), .A3(new_n462_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n653_));
  AND3_X1   g452(.A1(new_n652_), .A2(G22gat), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n652_), .B2(G22gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(G1327gat));
  NAND2_X1  g455(.A1(new_n628_), .A2(new_n587_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n567_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n467_), .A3(new_n508_), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n659_), .A2(G29gat), .A3(new_n463_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n618_), .A2(new_n587_), .A3(new_n620_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n608_), .A2(new_n610_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n467_), .B2(new_n664_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT43), .B(new_n663_), .C1(new_n438_), .C2(new_n466_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n661_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n370_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n671_), .B2(G29gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n660_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT109), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n677_), .B(new_n660_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n669_), .A2(new_n634_), .A3(new_n670_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G36gat), .ZN(new_n681_));
  INV_X1    g480(.A(new_n634_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n658_), .A2(new_n467_), .A3(new_n508_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n681_), .A2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT111), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n686_), .B1(new_n680_), .B2(G36gat), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n689_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n692_), .A2(new_n695_), .A3(KEYINPUT46), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n692_), .B2(KEYINPUT46), .ZN(new_n697_));
  OAI22_X1  g496(.A1(new_n691_), .A2(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(G1329gat));
  NAND4_X1  g497(.A1(new_n669_), .A2(G43gat), .A3(new_n643_), .A4(new_n670_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n331_), .B1(new_n659_), .B2(new_n334_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g501(.A1(new_n669_), .A2(new_n462_), .A3(new_n670_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G50gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n281_), .A2(G50gat), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT113), .Z(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n659_), .B2(new_n706_), .ZN(G1331gat));
  NOR2_X1   g506(.A1(new_n568_), .A2(new_n587_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n663_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT114), .Z(new_n710_));
  NOR2_X1   g509(.A1(new_n625_), .A2(new_n508_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n370_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n508_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n629_), .A2(new_n715_), .A3(new_n708_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(G57gat), .A3(new_n370_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(KEYINPUT115), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(KEYINPUT115), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n714_), .A2(new_n718_), .A3(new_n719_), .ZN(G1332gat));
  OR3_X1    g519(.A1(new_n712_), .A2(G64gat), .A3(new_n682_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n634_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G64gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(KEYINPUT48), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(KEYINPUT48), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(G1333gat));
  NAND2_X1  g525(.A1(new_n716_), .A2(new_n643_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G71gat), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT49), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT49), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n334_), .A2(G71gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT116), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n729_), .A2(new_n730_), .B1(new_n712_), .B2(new_n732_), .ZN(G1334gat));
  OR3_X1    g532(.A1(new_n712_), .A2(G78gat), .A3(new_n281_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n716_), .A2(new_n462_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G78gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(KEYINPUT50), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n736_), .A2(KEYINPUT50), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n657_), .A2(new_n568_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n711_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G85gat), .B1(new_n742_), .B2(new_n370_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n567_), .A2(new_n715_), .A3(new_n587_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n625_), .B2(new_n663_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n467_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n370_), .A2(G85gat), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT117), .Z(new_n749_));
  AOI21_X1  g548(.A(new_n743_), .B1(new_n747_), .B2(new_n749_), .ZN(G1336gat));
  INV_X1    g549(.A(G92gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n742_), .A2(new_n751_), .A3(new_n634_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n747_), .A2(new_n634_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n751_), .ZN(G1337gat));
  AOI21_X1  g553(.A(new_n532_), .B1(new_n747_), .B2(new_n643_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n742_), .A2(new_n643_), .A3(new_n543_), .ZN(new_n756_));
  OAI22_X1  g555(.A1(new_n755_), .A2(new_n756_), .B1(KEYINPUT118), .B2(KEYINPUT51), .ZN(new_n757_));
  NAND2_X1  g556(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1338gat));
  INV_X1    g558(.A(new_n744_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n462_), .B(new_n760_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762_));
  OAI21_X1  g561(.A(G106gat), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT119), .B1(new_n747_), .B2(new_n462_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n747_), .A2(KEYINPUT119), .A3(new_n462_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n762_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .A4(G106gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n742_), .A2(new_n533_), .A3(new_n462_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n774_), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  NAND4_X1  g575(.A1(new_n611_), .A2(new_n715_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n561_), .A2(new_n562_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n490_), .A2(new_n496_), .A3(new_n492_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n471_), .B1(new_n495_), .B2(new_n491_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT121), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n471_), .B2(new_n504_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n780_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n558_), .A2(new_n513_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n551_), .A2(new_n514_), .A3(new_n553_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(KEYINPUT55), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n560_), .B1(new_n554_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n786_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n786_), .A2(KEYINPUT58), .A3(new_n796_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n664_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n563_), .A2(new_n785_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n789_), .A2(new_n791_), .A3(new_n803_), .A4(KEYINPUT56), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n508_), .A2(new_n780_), .A3(new_n804_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n794_), .A2(KEYINPUT120), .A3(new_n795_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(new_n628_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n801_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n779_), .B1(new_n812_), .B2(new_n587_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n624_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n643_), .A2(new_n370_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n508_), .A2(new_n820_), .A3(G113gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n820_), .B2(G113gat), .ZN(new_n822_));
  INV_X1    g621(.A(new_n816_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n812_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n801_), .B(KEYINPUT122), .C1(new_n810_), .C2(new_n811_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n587_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n779_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n819_), .B(new_n822_), .C1(new_n829_), .C2(new_n817_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n829_), .B2(new_n508_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1340gat));
  OAI21_X1  g632(.A(new_n567_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n827_), .A2(new_n828_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n816_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(KEYINPUT59), .ZN(new_n837_));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  AND2_X1   g637(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n567_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT124), .B1(new_n829_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n619_), .B1(new_n812_), .B2(new_n824_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n779_), .B1(new_n844_), .B2(new_n826_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  NOR4_X1   g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n823_), .A4(new_n841_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n837_), .A2(new_n838_), .B1(new_n843_), .B2(new_n847_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n836_), .B2(new_n587_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n587_), .A2(new_n849_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n819_), .B(new_n851_), .C1(new_n829_), .C2(new_n817_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1342gat));
  INV_X1    g652(.A(G134gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n836_), .B2(new_n809_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n663_), .A2(new_n854_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n819_), .B(new_n856_), .C1(new_n829_), .C2(new_n817_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1343gat));
  NOR4_X1   g657(.A1(new_n634_), .A2(new_n463_), .A3(new_n281_), .A4(new_n643_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n835_), .A2(new_n508_), .A3(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g660(.A1(new_n835_), .A2(new_n567_), .A3(new_n859_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g662(.A1(new_n835_), .A2(new_n619_), .A3(new_n859_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  AND2_X1   g665(.A1(new_n835_), .A2(new_n859_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n664_), .A2(G162gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT125), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n835_), .A2(new_n628_), .A3(new_n859_), .ZN(new_n870_));
  INV_X1    g669(.A(G162gat), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n867_), .A2(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1347gat));
  NAND2_X1  g671(.A1(new_n634_), .A2(new_n371_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n462_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n813_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT126), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n813_), .B2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT22), .B(G169gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n508_), .A3(new_n881_), .ZN(new_n882_));
  AOI211_X1 g681(.A(KEYINPUT62), .B(new_n296_), .C1(new_n876_), .C2(new_n508_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n876_), .A2(new_n508_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(G169gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n882_), .B1(new_n883_), .B2(new_n886_), .ZN(G1348gat));
  INV_X1    g686(.A(new_n873_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(G176gat), .A3(new_n567_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n845_), .A2(new_n462_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n880_), .A2(new_n567_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n297_), .ZN(G1349gat));
  NOR2_X1   g691(.A1(new_n587_), .A2(new_n293_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n835_), .A2(new_n281_), .A3(new_n619_), .A4(new_n888_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n880_), .A2(new_n893_), .B1(new_n894_), .B2(new_n289_), .ZN(G1350gat));
  NOR2_X1   g694(.A1(new_n809_), .A2(new_n286_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n880_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n663_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n282_), .B2(new_n898_), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n682_), .A2(new_n464_), .A3(new_n643_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n835_), .A2(new_n900_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n901_), .A2(new_n207_), .A3(new_n715_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n900_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n845_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G197gat), .B1(new_n904_), .B2(new_n508_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n902_), .A2(new_n905_), .ZN(G1352gat));
  OAI21_X1  g705(.A(G204gat), .B1(new_n901_), .B2(new_n568_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n567_), .A2(new_n220_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT127), .B1(new_n904_), .B2(new_n908_), .ZN(new_n909_));
  AND4_X1   g708(.A1(KEYINPUT127), .A2(new_n835_), .A3(new_n900_), .A4(new_n908_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n907_), .B1(new_n909_), .B2(new_n910_), .ZN(G1353gat));
  XNOR2_X1  g710(.A(KEYINPUT63), .B(G211gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n901_), .A2(new_n587_), .A3(new_n912_), .ZN(new_n913_));
  OR2_X1    g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n904_), .B2(new_n619_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n901_), .B2(new_n663_), .ZN(new_n917_));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n904_), .A2(new_n918_), .A3(new_n628_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1355gat));
endmodule


