//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  INV_X1    g000(.A(G57gat), .ZN(new_n202_));
  INV_X1    g001(.A(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n210_), .A3(new_n205_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT11), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT12), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n217_), .A2(KEYINPUT69), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .A4(KEYINPUT68), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n224_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT7), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT6), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n219_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n234_), .B(new_n219_), .C1(new_n227_), .C2(new_n231_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT10), .B(G99gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(new_n236_), .B2(G106gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n229_), .A2(new_n230_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n221_), .A2(KEYINPUT10), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n221_), .A2(KEYINPUT10), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n239_), .B(new_n222_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n244_), .A2(new_n245_), .B1(G85gat), .B2(G92gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n217_), .B1(KEYINPUT66), .B2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(KEYINPUT66), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n243_), .B2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n222_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n231_), .B1(new_n252_), .B2(KEYINPUT64), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  INV_X1    g053(.A(new_n245_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n218_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n247_), .A2(KEYINPUT66), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n247_), .A2(KEYINPUT66), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n217_), .A4(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n253_), .A2(new_n254_), .A3(new_n260_), .A4(new_n242_), .ZN(new_n261_));
  AOI221_X4 g060(.A(KEYINPUT70), .B1(new_n233_), .B2(new_n235_), .C1(new_n251_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n233_), .A2(new_n235_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n216_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n251_), .A2(new_n261_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n214_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n215_), .B1(new_n269_), .B2(new_n214_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n264_), .A2(new_n265_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n214_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n268_), .B1(new_n276_), .B2(new_n270_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G120gat), .B(G148gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G204gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G176gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n273_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n282_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT71), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(KEYINPUT71), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n285_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n283_), .B(new_n284_), .C1(KEYINPUT71), .C2(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n292_));
  XOR2_X1   g091(.A(G15gat), .B(G22gat), .Z(new_n293_));
  XOR2_X1   g092(.A(KEYINPUT75), .B(G1gat), .Z(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G8gat), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n293_), .B1(new_n295_), .B2(KEYINPUT14), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n296_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G29gat), .B(G36gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n292_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n296_), .B(new_n297_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(KEYINPUT80), .A3(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G229gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n302_), .B(KEYINPUT15), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT81), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n307_), .A2(new_n313_), .A3(new_n308_), .A4(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n299_), .A2(new_n303_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(new_n314_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G141gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G169gat), .B(G197gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n311_), .A2(KEYINPUT81), .B1(new_n316_), .B2(new_n317_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT82), .A3(new_n314_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n324_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n312_), .A2(new_n318_), .A3(new_n314_), .A4(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT83), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n325_), .A2(new_n331_), .A3(new_n314_), .A4(new_n328_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n291_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  INV_X1    g135(.A(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT89), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT90), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT3), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n353_), .A2(new_n355_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n350_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n352_), .A2(new_n356_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n348_), .B(KEYINPUT1), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(new_n347_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n344_), .A2(KEYINPUT89), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n345_), .A2(new_n365_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n345_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n347_), .A2(new_n363_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n370_), .A2(new_n362_), .B1(new_n350_), .B2(new_n360_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n344_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(KEYINPUT102), .B(new_n368_), .C1(new_n373_), .C2(new_n366_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT102), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n372_), .A3(new_n375_), .A4(KEYINPUT4), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n341_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n341_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n340_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n369_), .A2(new_n372_), .A3(KEYINPUT4), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n368_), .A2(KEYINPUT102), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n376_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n378_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n379_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n340_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n380_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390_));
  XOR2_X1   g189(.A(G64gat), .B(G92gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(G211gat), .ZN(new_n398_));
  INV_X1    g197(.A(G218gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G211gat), .A2(G218gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT95), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT95), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n404_), .A3(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G197gat), .B(G204gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT21), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n408_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n406_), .A2(KEYINPUT96), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n407_), .A2(new_n408_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n407_), .B(KEYINPUT21), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT96), .B1(new_n415_), .B2(new_n406_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT24), .ZN(new_n418_));
  INV_X1    g217(.A(G169gat), .ZN(new_n419_));
  INV_X1    g218(.A(G176gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(KEYINPUT84), .A2(G183gat), .A3(G190gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT23), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n422_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n425_), .A2(new_n422_), .A3(new_n428_), .A4(new_n426_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n423_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n421_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT86), .B(new_n421_), .C1(new_n429_), .C2(new_n432_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT25), .B(G183gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT26), .B(G190gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n418_), .B1(G169gat), .B2(G176gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n419_), .A2(new_n420_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n437_), .A2(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT22), .B(G169gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n420_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G169gat), .A2(G176gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n423_), .A2(KEYINPUT23), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(G183gat), .A2(G190gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n446_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n417_), .B1(new_n442_), .B2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT103), .B(KEYINPUT20), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n415_), .A2(new_n406_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n421_), .A3(new_n441_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n413_), .A3(new_n411_), .A4(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n451_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n446_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n455_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n397_), .B1(new_n454_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n437_), .A2(new_n438_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n439_), .A2(new_n440_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n421_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n425_), .A2(new_n426_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n447_), .B1(new_n471_), .B2(KEYINPUT23), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT99), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT99), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n449_), .A2(new_n441_), .A3(new_n474_), .A4(new_n421_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n463_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n458_), .A2(new_n413_), .A3(new_n411_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n467_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n442_), .A2(new_n417_), .A3(new_n453_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n397_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n395_), .B1(new_n466_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n397_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n397_), .A2(new_n467_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n486_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT100), .B1(new_n454_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n486_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n473_), .A2(new_n475_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(new_n417_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT100), .ZN(new_n492_));
  INV_X1    g291(.A(new_n441_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n452_), .B1(new_n494_), .B2(new_n436_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n491_), .B(new_n492_), .C1(new_n417_), .C2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n485_), .A2(new_n488_), .A3(new_n395_), .A4(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n483_), .B1(new_n497_), .B2(KEYINPUT104), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n454_), .A2(new_n487_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n499_), .A2(new_n492_), .B1(new_n484_), .B2(new_n397_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT104), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n395_), .A4(new_n488_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n390_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n485_), .A2(new_n488_), .A3(new_n496_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n395_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(new_n390_), .A3(new_n497_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n389_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G71gat), .B(G99gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G15gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G227gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT87), .B(G43gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n442_), .A2(new_n453_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT30), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n495_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n519_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n516_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n345_), .A2(new_n367_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT31), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n525_), .B(new_n528_), .C1(new_n524_), .C2(new_n516_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n518_), .A2(new_n521_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT88), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n515_), .B1(new_n531_), .B2(new_n522_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n524_), .A2(new_n516_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n527_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT97), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(G228gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(G228gat), .ZN(new_n540_));
  AND2_X1   g339(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n541_));
  NOR2_X1   g340(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n539_), .B(new_n540_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n365_), .A2(KEYINPUT29), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n478_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n478_), .A2(new_n544_), .A3(new_n543_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n537_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n549_), .A2(new_n545_), .A3(new_n536_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n365_), .B2(KEYINPUT29), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n371_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G22gat), .B(G50gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n553_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT92), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(KEYINPUT92), .A3(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n549_), .A2(new_n545_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n566_), .A2(new_n537_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT98), .B1(new_n549_), .B2(new_n545_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n546_), .A2(new_n569_), .A3(new_n547_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n570_), .A3(new_n535_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n551_), .A2(new_n565_), .B1(new_n567_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n529_), .A2(new_n534_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT105), .B1(new_n509_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n497_), .A2(KEYINPUT104), .ZN(new_n575_));
  INV_X1    g374(.A(new_n483_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n502_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT27), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n507_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n529_), .A2(new_n534_), .A3(new_n572_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT105), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n389_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n574_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n571_), .A2(new_n567_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n564_), .ZN(new_n585_));
  OAI22_X1  g384(.A1(new_n585_), .A2(new_n562_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n509_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n466_), .A2(new_n482_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n395_), .A2(KEYINPUT32), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n380_), .A2(new_n387_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n504_), .A2(new_n590_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n587_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n340_), .B1(new_n373_), .B2(new_n341_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n383_), .B2(new_n341_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n387_), .B2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n384_), .A2(KEYINPUT33), .A3(new_n385_), .A4(new_n386_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n597_), .A2(new_n497_), .A3(new_n506_), .A4(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n593_), .A2(new_n599_), .B1(new_n534_), .B2(new_n529_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n588_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n335_), .B1(new_n583_), .B2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n309_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT34), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT35), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(KEYINPUT35), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n269_), .B2(new_n302_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n603_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n606_), .B1(new_n603_), .B2(new_n608_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT74), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G134gat), .B(G162gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(KEYINPUT36), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n611_), .B(new_n618_), .C1(KEYINPUT36), .C2(new_n616_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n616_), .A2(KEYINPUT36), .ZN(new_n620_));
  OAI221_X1 g419(.A(KEYINPUT74), .B1(new_n617_), .B2(new_n620_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(KEYINPUT37), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n214_), .B(KEYINPUT76), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n305_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n628_), .A2(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n629_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n299_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT77), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT77), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(new_n398_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT16), .B(G183gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n636_), .A2(KEYINPUT17), .A3(new_n637_), .A4(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n641_), .B(KEYINPUT17), .Z(new_n643_));
  AND3_X1   g442(.A1(new_n631_), .A2(KEYINPUT78), .A3(new_n634_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT78), .B1(new_n631_), .B2(new_n634_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT79), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT79), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n642_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n627_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n602_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n389_), .A2(new_n294_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(KEYINPUT38), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(KEYINPUT38), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n388_), .B1(new_n578_), .B2(new_n507_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n581_), .B1(new_n658_), .B2(new_n580_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n509_), .A2(KEYINPUT105), .A3(new_n573_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n601_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n335_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n642_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n649_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n622_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n663_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n389_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n656_), .A2(new_n657_), .A3(new_n671_), .ZN(G1324gat));
  INV_X1    g471(.A(G8gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n579_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n669_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT106), .B(KEYINPUT39), .Z(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n653_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n676_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1325gat));
  INV_X1    g481(.A(G15gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n529_), .A2(new_n534_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n669_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT41), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT41), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n653_), .A2(new_n683_), .A3(new_n685_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(G1326gat));
  INV_X1    g490(.A(G22gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n653_), .A2(new_n692_), .A3(new_n587_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n669_), .A2(new_n587_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G22gat), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT42), .B(new_n692_), .C1(new_n669_), .C2(new_n587_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(G1327gat));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n651_), .A2(new_n622_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n602_), .B2(new_n703_), .ZN(new_n704_));
  AOI22_X1  g503(.A1(new_n574_), .A2(new_n582_), .B1(new_n588_), .B2(new_n600_), .ZN(new_n705_));
  NOR4_X1   g504(.A1(new_n705_), .A2(KEYINPUT109), .A3(new_n335_), .A4(new_n702_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n388_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n661_), .A2(new_n709_), .A3(KEYINPUT43), .A4(new_n627_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n626_), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n705_), .B2(new_n626_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n710_), .A2(new_n712_), .A3(new_n662_), .A4(new_n651_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n715_), .A2(G29gat), .A3(new_n388_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n661_), .A2(new_n627_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n666_), .B1(new_n717_), .B2(new_n711_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n718_), .A2(KEYINPUT44), .A3(new_n662_), .A4(new_n710_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n708_), .B1(new_n716_), .B2(new_n719_), .ZN(G1328gat));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n579_), .A2(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n707_), .B2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n661_), .A2(new_n662_), .A3(new_n703_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT109), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n602_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n728_), .A2(new_n724_), .A3(new_n729_), .A4(new_n725_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n723_), .B1(new_n726_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(G36gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n579_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n719_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n721_), .A2(new_n722_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n732_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n736_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n719_), .A2(new_n715_), .A3(new_n674_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G36gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n728_), .A2(new_n729_), .A3(new_n725_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT45), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n742_), .A2(new_n730_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n738_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n737_), .A2(new_n744_), .ZN(G1329gat));
  NAND4_X1  g544(.A1(new_n719_), .A2(new_n715_), .A3(G43gat), .A4(new_n685_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n728_), .A2(new_n685_), .A3(new_n729_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(G43gat), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(KEYINPUT112), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT112), .B1(new_n747_), .B2(new_n748_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT47), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n746_), .B(new_n753_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1330gat));
  AOI21_X1  g554(.A(G50gat), .B1(new_n707_), .B2(new_n587_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n715_), .A2(G50gat), .A3(new_n587_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n705_), .A2(new_n291_), .A3(new_n334_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n652_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n388_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(new_n202_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n668_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n202_), .A2(KEYINPUT114), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n202_), .A2(KEYINPUT114), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n389_), .B(new_n765_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT113), .B(G57gat), .C1(new_n761_), .C2(new_n388_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n763_), .A2(new_n768_), .A3(new_n769_), .ZN(G1332gat));
  NAND3_X1  g569(.A1(new_n761_), .A2(new_n203_), .A3(new_n674_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G64gat), .B1(new_n765_), .B2(new_n579_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT48), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT48), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n765_), .B2(new_n684_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n778_), .ZN(new_n780_));
  INV_X1    g579(.A(G71gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n761_), .A2(new_n781_), .A3(new_n685_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n780_), .A3(new_n782_), .ZN(G1334gat));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n761_), .A2(new_n784_), .A3(new_n587_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G78gat), .B1(new_n765_), .B2(new_n572_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(KEYINPUT50), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(KEYINPUT50), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n785_), .B1(new_n787_), .B2(new_n788_), .ZN(G1335gat));
  AND2_X1   g588(.A1(new_n760_), .A2(new_n703_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n388_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT116), .Z(new_n792_));
  NOR2_X1   g591(.A1(new_n291_), .A2(new_n334_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n710_), .A2(new_n712_), .A3(new_n793_), .A4(new_n651_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n794_), .A2(new_n337_), .A3(new_n389_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n792_), .A2(new_n795_), .ZN(G1336gat));
  AOI21_X1  g595(.A(G92gat), .B1(new_n790_), .B2(new_n674_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n794_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n674_), .A2(G92gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(G1337gat));
  OAI211_X1 g599(.A(new_n790_), .B(new_n685_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G99gat), .B1(new_n794_), .B2(new_n684_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n790_), .A2(new_n222_), .A3(new_n587_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(G106gat), .C1(new_n794_), .C2(new_n572_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n718_), .A2(new_n587_), .A3(new_n710_), .A4(new_n793_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n806_), .B1(new_n809_), .B2(G106gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT53), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n805_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1339gat));
  NOR2_X1   g614(.A1(new_n674_), .A2(new_n389_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  INV_X1    g616(.A(new_n216_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n274_), .A2(KEYINPUT70), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n269_), .A2(new_n263_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n271_), .A2(new_n270_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n817_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n267_), .A2(KEYINPUT119), .A3(new_n270_), .A4(new_n271_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n268_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(KEYINPUT120), .A4(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n821_), .A2(new_n822_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(KEYINPUT121), .A3(KEYINPUT55), .A4(new_n268_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(KEYINPUT121), .A2(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(KEYINPUT121), .A2(KEYINPUT55), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n272_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n267_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n268_), .B1(new_n833_), .B2(new_n817_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT120), .B1(new_n834_), .B2(new_n824_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n282_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT56), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n282_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n837_), .A2(new_n283_), .A3(new_n334_), .A4(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n307_), .A2(new_n317_), .A3(new_n310_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n328_), .B1(new_n316_), .B2(new_n308_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n330_), .A2(new_n332_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n285_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT57), .B1(new_n845_), .B2(new_n667_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n847_), .B(new_n622_), .C1(new_n840_), .C2(new_n844_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n837_), .A2(new_n283_), .A3(new_n839_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(KEYINPUT58), .A4(new_n843_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n837_), .A2(new_n843_), .A3(new_n283_), .A4(new_n839_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT123), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n626_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n666_), .B1(new_n849_), .B2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n334_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n666_), .A2(new_n860_), .A3(new_n626_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n861_), .A2(new_n862_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n861_), .A2(KEYINPUT118), .A3(new_n862_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n580_), .B(new_n816_), .C1(new_n859_), .C2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT59), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n845_), .A2(new_n667_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n847_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n845_), .A2(new_n667_), .A3(KEYINPUT57), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n858_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n651_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n580_), .A4(new_n816_), .ZN(new_n879_));
  INV_X1    g678(.A(G113gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n334_), .B2(KEYINPUT124), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(KEYINPUT124), .B2(new_n880_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n870_), .A2(new_n879_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n334_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n880_), .B1(new_n869_), .B2(new_n884_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1340gat));
  INV_X1    g685(.A(new_n291_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n870_), .A2(new_n879_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G120gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n573_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n291_), .A2(KEYINPUT60), .ZN(new_n891_));
  MUX2_X1   g690(.A(new_n891_), .B(KEYINPUT60), .S(G120gat), .Z(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(new_n816_), .A3(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n893_), .ZN(G1341gat));
  NAND4_X1  g693(.A1(new_n870_), .A2(new_n879_), .A3(G127gat), .A4(new_n666_), .ZN(new_n895_));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n869_), .B2(new_n651_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1342gat));
  NAND4_X1  g697(.A1(new_n870_), .A2(new_n879_), .A3(G134gat), .A4(new_n627_), .ZN(new_n899_));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n869_), .B2(new_n667_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1343gat));
  NOR2_X1   g701(.A1(new_n685_), .A2(new_n572_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n877_), .A2(new_n816_), .A3(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT125), .B(G141gat), .ZN(new_n905_));
  OR3_X1    g704(.A1(new_n904_), .A2(new_n884_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n904_), .B2(new_n884_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1344gat));
  OR3_X1    g707(.A1(new_n904_), .A2(G148gat), .A3(new_n291_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G148gat), .B1(new_n904_), .B2(new_n291_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1345gat));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  INV_X1    g711(.A(new_n904_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n666_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n912_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n904_), .A2(new_n651_), .A3(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1346gat));
  INV_X1    g716(.A(G162gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n904_), .A2(new_n918_), .A3(new_n626_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n913_), .A2(new_n622_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n918_), .B2(new_n920_), .ZN(G1347gat));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n579_), .A2(new_n388_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n580_), .B(new_n923_), .C1(new_n859_), .C2(new_n868_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n922_), .B(G169gat), .C1(new_n924_), .C2(new_n884_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n877_), .A2(new_n334_), .A3(new_n580_), .A4(new_n923_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n922_), .B1(new_n927_), .B2(G169gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n334_), .A2(new_n443_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT126), .Z(new_n930_));
  OAI22_X1  g729(.A1(new_n926_), .A2(new_n928_), .B1(new_n924_), .B2(new_n930_), .ZN(G1348gat));
  NOR2_X1   g730(.A1(new_n924_), .A2(new_n291_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n420_), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n924_), .B2(new_n651_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n890_), .A2(new_n437_), .A3(new_n666_), .A4(new_n923_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n924_), .B2(new_n626_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n622_), .A2(new_n438_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n924_), .B2(new_n938_), .ZN(G1351gat));
  NAND3_X1  g738(.A1(new_n877_), .A2(new_n903_), .A3(new_n923_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941_), .B2(new_n334_), .ZN(new_n942_));
  INV_X1    g741(.A(G197gat), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n940_), .A2(new_n943_), .A3(new_n884_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n942_), .A2(new_n944_), .ZN(G1352gat));
  NAND2_X1  g744(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n941_), .A2(new_n887_), .A3(new_n946_), .ZN(new_n947_));
  OAI211_X1 g746(.A(KEYINPUT127), .B(G204gat), .C1(new_n940_), .C2(new_n291_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1353gat));
  XOR2_X1   g748(.A(KEYINPUT63), .B(G211gat), .Z(new_n950_));
  NAND3_X1  g749(.A1(new_n941_), .A2(new_n666_), .A3(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n940_), .B2(new_n651_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1354gat));
  NOR3_X1   g753(.A1(new_n940_), .A2(new_n399_), .A3(new_n626_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n941_), .A2(new_n622_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n399_), .B2(new_n956_), .ZN(G1355gat));
endmodule


