//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  XOR2_X1   g001(.A(G85gat), .B(G92gat), .Z(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n203_), .B1(new_n206_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT8), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT10), .B(G99gat), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  AOI22_X1  g012(.A1(KEYINPUT9), .A2(new_n203_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT9), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n209_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n211_), .A2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(G78gat), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  INV_X1    g023(.A(G71gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G78gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n223_), .B(new_n229_), .C1(KEYINPUT11), .C2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT67), .ZN(new_n232_));
  INV_X1    g031(.A(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G57gat), .ZN(new_n234_));
  INV_X1    g033(.A(G57gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G64gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT11), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n223_), .A4(new_n229_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n232_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n232_), .B2(new_n240_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n221_), .A2(new_n222_), .A3(G78gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(new_n237_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n239_), .B1(new_n248_), .B2(new_n223_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n231_), .A2(KEYINPUT67), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n241_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n232_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT68), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n220_), .B1(new_n246_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT69), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(KEYINPUT68), .A3(new_n252_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n245_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n211_), .A2(new_n219_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n256_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n220_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n255_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G230gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n251_), .A2(KEYINPUT70), .A3(new_n252_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n211_), .B2(new_n219_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n259_), .A2(new_n268_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n267_), .B1(new_n260_), .B2(new_n220_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n263_), .A2(new_n267_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G120gat), .B(G148gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G176gat), .B(G204gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n263_), .A2(new_n267_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n259_), .A2(new_n268_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n272_), .A2(new_n273_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n275_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n288_), .A3(new_n282_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(KEYINPUT13), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  INV_X1    g090(.A(G1gat), .ZN(new_n292_));
  INV_X1    g091(.A(G8gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G29gat), .B(G36gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n297_), .B(new_n300_), .Z(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(G229gat), .A3(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n300_), .B(KEYINPUT15), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n297_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n297_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n300_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT77), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G113gat), .B(G141gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(G169gat), .B(G197gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n310_), .A2(new_n313_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT13), .ZN(new_n318_));
  INV_X1    g117(.A(new_n289_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(new_n283_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n290_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT23), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(G183gat), .B2(G190gat), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  INV_X1    g124(.A(G169gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT79), .B1(new_n326_), .B2(KEYINPUT22), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT22), .B(G169gat), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n325_), .B(new_n327_), .C1(new_n328_), .C2(KEYINPUT79), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n323_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n326_), .A2(new_n325_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(KEYINPUT24), .A3(new_n330_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G190gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(KEYINPUT78), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT78), .B1(new_n343_), .B2(G190gat), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n331_), .B1(new_n339_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT81), .ZN(new_n348_));
  XOR2_X1   g147(.A(G71gat), .B(G99gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n346_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT80), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT30), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT31), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n351_), .A2(new_n355_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT82), .B1(new_n356_), .B2(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G127gat), .B(G134gat), .Z(new_n363_));
  XOR2_X1   g162(.A(G113gat), .B(G120gat), .Z(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n365_), .A3(new_n361_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G155gat), .B(G162gat), .Z(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT85), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n384_), .A2(KEYINPUT84), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT84), .B1(new_n384_), .B2(new_n385_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n374_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n379_), .B(new_n382_), .C1(new_n387_), .C2(new_n386_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT86), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n374_), .ZN(new_n393_));
  INV_X1    g192(.A(G155gat), .ZN(new_n394_));
  INV_X1    g193(.A(G162gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT1), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT1), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(G155gat), .A3(G162gat), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n396_), .B(new_n398_), .C1(G155gat), .C2(G162gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(G141gat), .B(G148gat), .Z(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(KEYINPUT83), .A3(new_n400_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n390_), .A2(new_n393_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT87), .B(G204gat), .ZN(new_n410_));
  INV_X1    g209(.A(G197gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G218gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G211gat), .ZN(new_n414_));
  INV_X1    g213(.A(G211gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G218gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT21), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT88), .B1(new_n412_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(G204gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT87), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G204gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n408_), .B1(new_n424_), .B2(G197gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT21), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n412_), .A2(new_n427_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n421_), .A2(new_n423_), .A3(new_n411_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(G197gat), .B2(G204gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n417_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n419_), .A2(new_n429_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n373_), .B1(new_n407_), .B2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G78gat), .B(G106gat), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n403_), .A2(new_n404_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n391_), .A2(new_n392_), .A3(new_n374_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n392_), .B1(new_n391_), .B2(new_n374_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT29), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n430_), .A2(new_n433_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n412_), .A2(new_n418_), .A3(KEYINPUT88), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n426_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT89), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n434_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n373_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n442_), .A2(new_n447_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n435_), .A2(new_n437_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n437_), .B1(new_n435_), .B2(new_n451_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT28), .B1(new_n441_), .B2(KEYINPUT29), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT28), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n405_), .A2(new_n456_), .A3(new_n406_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G22gat), .B(G50gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n455_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n461_));
  OAI22_X1  g260(.A1(new_n453_), .A2(new_n454_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n435_), .A2(new_n451_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n436_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n460_), .A2(new_n461_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n452_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G29gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G85gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n441_), .A2(new_n365_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n390_), .A2(new_n393_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n366_), .A3(new_n438_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n473_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n474_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n474_), .B2(KEYINPUT4), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n366_), .B1(new_n475_), .B2(new_n438_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n478_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n474_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT92), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n480_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT94), .B1(new_n490_), .B2(KEYINPUT33), .ZN(new_n491_));
  INV_X1    g290(.A(new_n480_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n487_), .A2(KEYINPUT92), .A3(new_n488_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT92), .B1(new_n487_), .B2(new_n488_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G8gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT18), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G226gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT19), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n342_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(G183gat), .ZN(new_n511_));
  INV_X1    g310(.A(G183gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT25), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT90), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n509_), .A2(new_n514_), .A3(new_n340_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n338_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(KEYINPUT91), .A3(new_n338_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n336_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n328_), .A2(new_n325_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n324_), .A2(new_n330_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n507_), .B1(new_n523_), .B2(new_n446_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n447_), .A2(new_n449_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n346_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n506_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n447_), .A2(new_n449_), .A3(new_n346_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n520_), .A2(new_n434_), .A3(new_n522_), .ZN(new_n530_));
  AND4_X1   g329(.A1(KEYINPUT20), .A2(new_n529_), .A3(new_n506_), .A4(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n503_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n522_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n335_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(new_n519_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT20), .B1(new_n535_), .B2(new_n434_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n346_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n505_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n507_), .B1(new_n535_), .B2(new_n434_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(new_n506_), .A3(new_n529_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n502_), .A3(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n474_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n478_), .B1(new_n474_), .B2(KEYINPUT4), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n472_), .B(new_n542_), .C1(new_n482_), .C2(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n532_), .A2(new_n541_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n490_), .A2(KEYINPUT33), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n491_), .A2(new_n498_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n477_), .A2(new_n479_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n495_), .B1(new_n549_), .B2(new_n473_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n502_), .A2(KEYINPUT32), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n528_), .A2(new_n531_), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n524_), .A2(new_n506_), .A3(new_n527_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n539_), .A2(new_n529_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(new_n506_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n467_), .B1(new_n547_), .B2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n493_), .A2(new_n494_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n472_), .B1(new_n559_), .B2(new_n548_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n467_), .A2(new_n495_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n503_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(KEYINPUT27), .A3(new_n541_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n532_), .A2(new_n541_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n370_), .B1(new_n558_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n567_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n550_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n467_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n570_), .A2(new_n369_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n321_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT36), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n258_), .A2(new_n303_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT34), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT35), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT72), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(KEYINPUT35), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n220_), .B2(new_n300_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n586_), .B1(new_n581_), .B2(new_n588_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n578_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n577_), .A2(KEYINPUT36), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n589_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n592_), .A2(new_n595_), .A3(new_n596_), .A4(KEYINPUT37), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  AND2_X1   g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n297_), .B(new_n610_), .ZN(new_n611_));
  AOI211_X1 g410(.A(new_n608_), .B(new_n609_), .C1(new_n611_), .C2(new_n260_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n260_), .A2(new_n611_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n272_), .A2(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n272_), .A2(new_n611_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n608_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT76), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n612_), .A2(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n601_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n574_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n571_), .A2(KEYINPUT96), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n571_), .A2(KEYINPUT96), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(new_n292_), .A3(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT97), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT97), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(KEYINPUT38), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n592_), .A2(new_n595_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n321_), .A2(new_n620_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G1gat), .B1(new_n638_), .B2(new_n571_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n633_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT38), .B1(new_n631_), .B2(new_n632_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n202_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(KEYINPUT98), .A3(new_n639_), .A4(new_n633_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n624_), .A2(new_n293_), .A3(new_n567_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n636_), .A2(new_n567_), .A3(new_n637_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  AND4_X1   g447(.A1(KEYINPUT99), .A2(new_n647_), .A3(new_n648_), .A4(G8gat), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n293_), .B1(new_n650_), .B2(KEYINPUT39), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n647_), .A2(new_n651_), .B1(KEYINPUT99), .B2(new_n648_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n646_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n638_), .B2(new_n370_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT41), .Z(new_n656_));
  INV_X1    g455(.A(G15gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n624_), .A2(new_n657_), .A3(new_n369_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n624_), .A2(new_n660_), .A3(new_n467_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G22gat), .B1(new_n638_), .B2(new_n572_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT42), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(KEYINPUT42), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT100), .ZN(G1327gat));
  NOR2_X1   g465(.A1(new_n634_), .A2(new_n621_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n574_), .A2(KEYINPUT102), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT102), .B1(new_n574_), .B2(new_n667_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n550_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n569_), .A2(new_n573_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n599_), .A2(new_n600_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n601_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n321_), .A2(new_n621_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  INV_X1    g482(.A(new_n681_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n683_), .B(new_n684_), .C1(new_n675_), .C2(new_n679_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n629_), .A2(G29gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n671_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  XNOR2_X1  g487(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(G36gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n686_), .B2(new_n567_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n570_), .A2(G36gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT104), .B1(new_n670_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n321_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n672_), .A2(new_n697_), .A3(new_n667_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n574_), .A2(KEYINPUT102), .A3(new_n667_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n695_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n694_), .B1(new_n696_), .B2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n670_), .A2(KEYINPUT104), .A3(new_n695_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n703_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n693_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n690_), .B1(new_n692_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n680_), .A2(new_n681_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n683_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n681_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n567_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G36gat), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n715_), .A2(new_n708_), .A3(new_n705_), .A4(new_n689_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n710_), .A2(new_n716_), .ZN(G1329gat));
  AND2_X1   g516(.A1(new_n369_), .A2(G43gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n700_), .A2(new_n369_), .A3(new_n701_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT106), .B(G43gat), .Z(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT107), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n719_), .A2(new_n723_), .A3(new_n720_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n686_), .A2(new_n718_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n670_), .B2(new_n467_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n467_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n686_), .B2(new_n729_), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n290_), .A2(new_n320_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n636_), .A2(new_n621_), .A3(new_n316_), .A4(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n732_), .A2(new_n235_), .A3(new_n571_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n731_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n317_), .B(new_n734_), .C1(new_n569_), .C2(new_n573_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n623_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n628_), .B1(new_n736_), .B2(KEYINPUT109), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(KEYINPUT109), .B2(new_n736_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n733_), .B1(new_n738_), .B2(new_n235_), .ZN(G1332gat));
  OAI21_X1  g538(.A(G64gat), .B1(new_n732_), .B2(new_n570_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n567_), .A2(new_n233_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n736_), .B2(new_n743_), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n732_), .B2(new_n370_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT49), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n369_), .A2(new_n225_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n736_), .B2(new_n747_), .ZN(G1334gat));
  OAI21_X1  g547(.A(G78gat), .B1(new_n732_), .B2(new_n572_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT50), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n467_), .A2(new_n227_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n736_), .B2(new_n751_), .ZN(G1335gat));
  NAND3_X1  g551(.A1(new_n731_), .A2(new_n620_), .A3(new_n316_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n680_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n571_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n735_), .A2(new_n667_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n215_), .A3(new_n629_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1336gat));
  OAI21_X1  g559(.A(G92gat), .B1(new_n755_), .B2(new_n570_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n567_), .A2(new_n216_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n757_), .B2(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT111), .Z(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n755_), .B2(new_n370_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n369_), .A2(new_n212_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n757_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT51), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n767_), .B(new_n769_), .Z(G1338gat));
  AOI21_X1  g569(.A(KEYINPUT43), .B1(new_n674_), .B2(KEYINPUT101), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n677_), .A2(new_n678_), .A3(new_n676_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n467_), .B(new_n754_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G106gat), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n572_), .B(new_n753_), .C1(new_n675_), .C2(new_n679_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT113), .B(new_n777_), .C1(new_n779_), .C2(new_n213_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n758_), .A2(new_n213_), .A3(new_n467_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT53), .B1(new_n778_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT113), .B1(new_n779_), .B2(new_n213_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(KEYINPUT52), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n780_), .A4(new_n781_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(new_n788_), .ZN(G1339gat));
  OAI21_X1  g588(.A(KEYINPUT114), .B1(new_n620_), .B2(new_n317_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n621_), .A2(new_n791_), .A3(new_n316_), .ZN(new_n792_));
  AND4_X1   g591(.A1(new_n599_), .A2(new_n790_), .A3(new_n600_), .A4(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n734_), .A3(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n599_), .A2(new_n600_), .A3(new_n792_), .A4(new_n790_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT54), .B1(new_n796_), .B2(new_n731_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  INV_X1    g598(.A(new_n308_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n304_), .A2(new_n306_), .A3(new_n800_), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n313_), .B(new_n801_), .C1(new_n301_), .C2(new_n308_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n314_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n284_), .B2(new_n289_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n274_), .A2(new_n255_), .A3(new_n262_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n267_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n274_), .A2(KEYINPUT55), .A3(new_n275_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n288_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n808_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n281_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n281_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n811_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n281_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n316_), .B1(new_n276_), .B2(new_n282_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n805_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n799_), .B1(new_n821_), .B2(new_n635_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n819_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n806_), .A2(new_n267_), .B1(new_n288_), .B2(new_n809_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n813_), .B(new_n282_), .C1(new_n824_), .C2(new_n808_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n281_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n823_), .B1(new_n827_), .B2(new_n815_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT57), .B(new_n634_), .C1(new_n828_), .C2(new_n805_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n319_), .B2(new_n804_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n289_), .A2(new_n803_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n834_), .B2(new_n827_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n814_), .A2(new_n816_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT58), .A3(new_n833_), .A4(new_n831_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n837_), .A3(new_n673_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n822_), .A2(new_n829_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n621_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n822_), .A2(new_n829_), .A3(KEYINPUT117), .A4(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n798_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n570_), .A2(new_n572_), .A3(new_n369_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n628_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n317_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n839_), .A2(new_n620_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n798_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n845_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n317_), .B(new_n854_), .C1(new_n847_), .C2(new_n853_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n849_), .B1(new_n856_), .B2(new_n848_), .ZN(G1340gat));
  OAI211_X1 g656(.A(new_n731_), .B(new_n854_), .C1(new_n847_), .C2(new_n853_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT118), .B(G120gat), .Z(new_n860_));
  INV_X1    g659(.A(new_n847_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n734_), .B2(KEYINPUT60), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(KEYINPUT60), .B2(new_n860_), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n859_), .A2(new_n860_), .B1(new_n861_), .B2(new_n863_), .ZN(G1341gat));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n847_), .A2(new_n865_), .A3(new_n621_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n621_), .B(new_n854_), .C1(new_n847_), .C2(new_n853_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n868_), .B2(new_n865_), .ZN(G1342gat));
  INV_X1    g668(.A(G134gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n847_), .A2(new_n870_), .A3(new_n635_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n673_), .B(new_n854_), .C1(new_n847_), .C2(new_n853_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n870_), .ZN(G1343gat));
  NAND4_X1  g673(.A1(new_n629_), .A2(new_n467_), .A3(new_n570_), .A4(new_n370_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n839_), .A2(new_n840_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n620_), .A3(new_n842_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n851_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n317_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n731_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n878_), .B2(new_n621_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n843_), .A2(KEYINPUT119), .A3(new_n620_), .A4(new_n875_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n877_), .A2(new_n851_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n875_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n621_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT119), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n878_), .A2(new_n885_), .A3(new_n621_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n883_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n888_), .A2(new_n894_), .ZN(G1346gat));
  INV_X1    g694(.A(new_n878_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G162gat), .B1(new_n896_), .B2(new_n601_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n878_), .A2(new_n395_), .A3(new_n635_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n798_), .B1(new_n620_), .B2(new_n839_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n370_), .A2(new_n570_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n628_), .A2(new_n572_), .A3(new_n902_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n901_), .A2(new_n316_), .A3(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n900_), .B1(new_n904_), .B2(new_n326_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n903_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n852_), .A2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT62), .B(G169gat), .C1(new_n907_), .C2(new_n316_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n328_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n905_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n905_), .A2(new_n908_), .A3(KEYINPUT120), .A4(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n901_), .A2(new_n903_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G176gat), .B1(new_n915_), .B2(new_n731_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n843_), .A2(new_n903_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n734_), .A2(new_n325_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(KEYINPUT121), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n921_), .A3(new_n918_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n916_), .B1(new_n920_), .B2(new_n922_), .ZN(G1349gat));
  AOI21_X1  g722(.A(new_n620_), .B1(new_n514_), .B2(new_n509_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n915_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G183gat), .B1(new_n917_), .B2(new_n621_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n907_), .B2(new_n601_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n915_), .A2(new_n635_), .A3(new_n340_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1351gat));
  OR2_X1    g731(.A1(new_n561_), .A2(new_n369_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n933_), .A2(KEYINPUT123), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(KEYINPUT123), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n934_), .A2(new_n567_), .A3(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n843_), .A2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n317_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT124), .B(G197gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1352gat));
  NAND2_X1  g739(.A1(new_n937_), .A2(new_n731_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n410_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n420_), .B2(new_n941_), .ZN(G1353gat));
  NAND2_X1  g742(.A1(new_n937_), .A2(new_n621_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT63), .B(G211gat), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n944_), .B2(new_n947_), .ZN(G1354gat));
  NOR3_X1   g747(.A1(new_n843_), .A2(new_n634_), .A3(new_n936_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(KEYINPUT125), .B(G218gat), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n936_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n673_), .A2(new_n950_), .ZN(new_n953_));
  XOR2_X1   g752(.A(new_n953_), .B(KEYINPUT126), .Z(new_n954_));
  AND3_X1   g753(.A1(new_n889_), .A2(new_n952_), .A3(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(KEYINPUT127), .B1(new_n951_), .B2(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n937_), .A2(new_n954_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n957_), .B(new_n958_), .C1(new_n949_), .C2(new_n950_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n956_), .A2(new_n959_), .ZN(G1355gat));
endmodule


