//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_;
  INV_X1    g000(.A(G155gat), .ZN(new_n202_));
  INV_X1    g001(.A(G162gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT82), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT82), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT87), .A4(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  INV_X1    g013(.A(G141gat), .ZN(new_n215_));
  INV_X1    g014(.A(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  OAI22_X1  g016(.A1(KEYINPUT85), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n222_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n219_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT88), .B1(new_n212_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n225_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n229_), .A2(KEYINPUT2), .B1(KEYINPUT85), .B2(KEYINPUT3), .ZN(new_n230_));
  INV_X1    g029(.A(new_n226_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n218_), .A4(new_n217_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT88), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G141gat), .B(G148gat), .Z(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT83), .B1(new_n207_), .B2(KEYINPUT1), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT83), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(G155gat), .A4(G162gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n204_), .A2(new_n241_), .A3(new_n206_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n235_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT84), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  OAI211_X1 g044(.A(KEYINPUT84), .B(new_n235_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n228_), .A2(new_n234_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G22gat), .B(G50gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT28), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n249_), .B(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n228_), .A2(new_n234_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n246_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT92), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(KEYINPUT29), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT92), .B1(new_n247_), .B2(new_n248_), .ZN(new_n258_));
  INV_X1    g057(.A(G197gat), .ZN(new_n259_));
  AND2_X1   g058(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G197gat), .A2(G204gat), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n262_), .A2(KEYINPUT21), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G211gat), .B(G218gat), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT89), .B(G204gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(G197gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT90), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(G197gat), .B1(new_n260_), .B2(new_n261_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n274_), .A2(KEYINPUT90), .A3(new_n272_), .A4(new_n268_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n265_), .B(new_n267_), .C1(new_n273_), .C2(new_n276_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n271_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n257_), .A2(new_n258_), .A3(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(G228gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT91), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n277_), .A2(KEYINPUT91), .A3(new_n279_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n282_), .B1(new_n255_), .B2(KEYINPUT29), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n281_), .A2(new_n282_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G78gat), .B(G106gat), .Z(new_n289_));
  OAI21_X1  g088(.A(new_n252_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n281_), .A2(new_n282_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n289_), .B(KEYINPUT93), .Z(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n287_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT94), .B1(new_n290_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n293_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n289_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n288_), .A2(new_n292_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .A4(new_n252_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n252_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n292_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n294_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT26), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n306_), .A2(KEYINPUT26), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT80), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G183gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT79), .B1(new_n311_), .B2(KEYINPUT25), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(new_n307_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT25), .B(G183gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n310_), .B(new_n314_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT23), .ZN(new_n319_));
  INV_X1    g118(.A(G169gat), .ZN(new_n320_));
  INV_X1    g119(.A(G176gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n321_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT24), .A3(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n324_), .A2(KEYINPUT24), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n317_), .A2(new_n319_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT30), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n319_), .B1(G183gat), .B2(G190gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G169gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n322_), .B1(new_n330_), .B2(new_n321_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n327_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n328_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n334_));
  OAI21_X1  g133(.A(G43gat), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n327_), .A2(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT30), .ZN(new_n337_));
  INV_X1    g136(.A(G43gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n327_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G15gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  AND3_X1   g143(.A1(new_n335_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT81), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n335_), .A2(new_n340_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n344_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n335_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  INV_X1    g153(.A(G113gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G120gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT31), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n347_), .A2(new_n353_), .A3(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT81), .B(new_n359_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n305_), .A2(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n361_), .A2(new_n362_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n365_), .A2(new_n304_), .A3(new_n295_), .A4(new_n301_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n247_), .A2(new_n358_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n247_), .A2(new_n358_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(KEYINPUT99), .A2(new_n370_), .B1(new_n371_), .B2(KEYINPUT4), .ZN(new_n372_));
  INV_X1    g171(.A(new_n358_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n255_), .A2(KEYINPUT99), .A3(new_n373_), .A4(KEYINPUT4), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n369_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n255_), .A2(new_n373_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n377_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G85gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(G1gat), .B(G29gat), .Z(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n376_), .A2(new_n379_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n255_), .A2(KEYINPUT99), .A3(new_n373_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n247_), .B2(new_n358_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n374_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n378_), .B1(new_n390_), .B2(new_n369_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(new_n384_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n386_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT27), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT18), .B(G64gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G92gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n396_), .B(new_n397_), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n277_), .A2(KEYINPUT91), .A3(new_n279_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT91), .B1(new_n277_), .B2(new_n279_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n336_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n331_), .B(KEYINPUT97), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n329_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT26), .B(G190gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT95), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n316_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n323_), .A2(new_n324_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n407_), .A2(new_n319_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n404_), .A2(new_n412_), .A3(new_n277_), .A4(new_n279_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT19), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n284_), .A2(new_n285_), .A3(new_n332_), .A4(new_n327_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n404_), .A2(new_n412_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n280_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n419_), .A2(KEYINPUT20), .A3(new_n416_), .A4(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n399_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n286_), .B2(new_n336_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(KEYINPUT20), .A3(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n417_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n398_), .B(KEYINPUT101), .Z(new_n430_));
  AOI211_X1 g229(.A(new_n394_), .B(new_n423_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n416_), .B1(new_n425_), .B2(new_n413_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n422_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n398_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n418_), .A2(new_n422_), .A3(new_n399_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT27), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n367_), .A2(new_n393_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n429_), .A2(KEYINPUT32), .A3(new_n398_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n398_), .A2(KEYINPUT32), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n439_), .B(new_n441_), .C1(new_n392_), .C2(new_n386_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT98), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n418_), .A2(new_n422_), .A3(new_n399_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n423_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n434_), .A2(new_n435_), .A3(KEYINPUT98), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n376_), .A2(KEYINPUT33), .A3(new_n379_), .A4(new_n384_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n390_), .A2(new_n368_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n377_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n383_), .A3(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n385_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT100), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT100), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n385_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n442_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n305_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n363_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n438_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G230gat), .A2(G233gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT64), .Z(new_n464_));
  NAND2_X1  g263(.A1(G57gat), .A2(G64gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G57gat), .A2(G64gat), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT68), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n469_));
  INV_X1    g268(.A(G57gat), .ZN(new_n470_));
  INV_X1    g269(.A(G64gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n472_), .B2(new_n465_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT11), .B1(new_n468_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G71gat), .B(G78gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT68), .B1(new_n466_), .B2(new_n467_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT11), .B(new_n475_), .C1(new_n468_), .C2(new_n473_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT10), .B(G99gat), .Z(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G85gat), .B(G92gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT9), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n490_));
  NOR2_X1   g289(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(G92gat), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AND3_X1   g291(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n486_), .A2(new_n488_), .A3(new_n492_), .A4(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  INV_X1    g296(.A(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(new_n485_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT7), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n497_), .A2(new_n501_), .A3(new_n498_), .A4(new_n485_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n495_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n487_), .A3(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n503_), .A2(new_n487_), .A3(new_n508_), .A4(new_n504_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n483_), .A2(new_n496_), .A3(new_n507_), .A4(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT69), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n481_), .A2(new_n482_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n507_), .A2(new_n496_), .A3(new_n509_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n511_), .A2(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT69), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n510_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT70), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n464_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n464_), .B1(new_n514_), .B2(new_n513_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT72), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n513_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n481_), .A2(KEYINPUT71), .A3(new_n482_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT71), .B1(new_n481_), .B2(new_n482_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT12), .B(new_n514_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n521_), .A2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G120gat), .B(G148gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G176gat), .B(G204gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n519_), .A2(new_n529_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n519_), .B2(new_n529_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT13), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(KEYINPUT13), .A3(new_n538_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G29gat), .B(G36gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n338_), .ZN(new_n544_));
  INV_X1    g343(.A(G50gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT15), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n544_), .B(G50gat), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552_));
  INV_X1    g351(.A(G1gat), .ZN(new_n553_));
  INV_X1    g352(.A(G8gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G1gat), .B(G8gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n548_), .A2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n548_), .B(new_n558_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n565_), .A2(new_n563_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n320_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n259_), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n564_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT78), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT78), .B(new_n569_), .C1(new_n564_), .C2(new_n566_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n542_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n462_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT74), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT74), .B1(new_n580_), .B2(new_n581_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n551_), .A2(new_n514_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n514_), .A2(new_n548_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n580_), .A2(new_n581_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n584_), .B(new_n585_), .C1(new_n586_), .C2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n551_), .A2(new_n514_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n591_), .A2(new_n583_), .A3(new_n582_), .A4(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT76), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT75), .B(G190gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G218gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(G134gat), .B(G162gat), .Z(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n600_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n594_), .A2(KEYINPUT76), .A3(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n590_), .A2(KEYINPUT36), .A3(new_n599_), .A4(new_n593_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT37), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n602_), .B1(new_n594_), .B2(KEYINPUT76), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n608_), .B(new_n600_), .C1(new_n590_), .C2(new_n593_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT37), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n604_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n558_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n483_), .ZN(new_n615_));
  XOR2_X1   g414(.A(G127gat), .B(G155gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G183gat), .B(G211gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n615_), .B1(KEYINPUT17), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(KEYINPUT71), .A3(KEYINPUT17), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n606_), .A2(new_n612_), .A3(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n577_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n393_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n553_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT102), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n628_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT104), .ZN(new_n632_));
  INV_X1    g431(.A(new_n623_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n577_), .A2(new_n633_), .A3(new_n605_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT103), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(new_n626_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n630_), .B(new_n632_), .C1(new_n553_), .C2(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(new_n437_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n625_), .A2(new_n554_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n634_), .A2(new_n638_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G8gat), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT39), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(KEYINPUT39), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n635_), .B2(new_n365_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT41), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n625_), .A2(new_n646_), .A3(new_n365_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT105), .Z(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n635_), .B2(new_n305_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT42), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n625_), .A2(new_n652_), .A3(new_n305_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(new_n577_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n605_), .A2(new_n633_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT108), .Z(new_n659_));
  AND2_X1   g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(G29gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n626_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n606_), .A2(new_n612_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n606_), .A2(new_n612_), .A3(KEYINPUT106), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n663_), .B1(new_n462_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n611_), .B1(new_n610_), .B2(new_n604_), .ZN(new_n670_));
  AND4_X1   g469(.A1(new_n611_), .A2(new_n601_), .A3(new_n603_), .A4(new_n604_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT43), .B(new_n672_), .C1(new_n438_), .C2(new_n461_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n576_), .B(new_n633_), .C1(new_n669_), .C2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT107), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n393_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n662_), .B1(new_n679_), .B2(new_n661_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT109), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n683_));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n660_), .A2(new_n683_), .A3(new_n684_), .A4(new_n638_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n657_), .A2(new_n684_), .A3(new_n638_), .A4(new_n659_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT45), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n437_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n682_), .B(new_n688_), .C1(new_n689_), .C2(new_n684_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n681_), .A2(KEYINPUT109), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n691_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n685_), .A2(new_n687_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n674_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT44), .B1(new_n674_), .B2(KEYINPUT107), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n638_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n697_), .B2(G36gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n693_), .B1(new_n698_), .B2(new_n682_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n692_), .A2(new_n699_), .ZN(G1329gat));
  OAI21_X1  g499(.A(new_n365_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n363_), .A2(G43gat), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n701_), .A2(G43gat), .B1(new_n660_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g503(.A1(new_n660_), .A2(new_n545_), .A3(new_n305_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n305_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G50gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1331gat));
  INV_X1    g509(.A(new_n541_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n539_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n575_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n462_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n605_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(new_n623_), .A3(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(G57gat), .A3(new_n626_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT111), .Z(new_n719_));
  INV_X1    g518(.A(new_n624_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n715_), .A2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n470_), .B1(new_n721_), .B2(new_n393_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n719_), .A2(KEYINPUT112), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1332gat));
  AOI21_X1  g526(.A(new_n471_), .B1(new_n717_), .B2(new_n638_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT48), .Z(new_n729_));
  INV_X1    g528(.A(new_n721_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n471_), .A3(new_n638_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n717_), .B2(new_n365_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT49), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n733_), .A3(new_n365_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1334gat));
  INV_X1    g536(.A(G78gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n717_), .B2(new_n305_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT50), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n738_), .A3(new_n305_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  AND2_X1   g541(.A1(new_n715_), .A2(new_n659_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n626_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n714_), .A2(new_n633_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT113), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(new_n747_), .C1(new_n669_), .C2(new_n673_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n745_), .B(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n669_), .A2(new_n673_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT114), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n748_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n491_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n393_), .B1(new_n754_), .B2(new_n489_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n744_), .B1(new_n753_), .B2(new_n755_), .ZN(G1336gat));
  AOI21_X1  g555(.A(G92gat), .B1(new_n743_), .B2(new_n638_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n638_), .A2(G92gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n753_), .B2(new_n758_), .ZN(G1337gat));
  NAND3_X1  g558(.A1(new_n748_), .A2(new_n752_), .A3(new_n365_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G99gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n743_), .A2(new_n484_), .A3(new_n365_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n743_), .A2(new_n485_), .A3(new_n305_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n750_), .A2(new_n751_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n305_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n768_), .B2(G106gat), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT52), .B(new_n485_), .C1(new_n767_), .C2(new_n305_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n765_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n765_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  INV_X1    g574(.A(new_n366_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n638_), .A2(new_n393_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n464_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n517_), .B2(new_n528_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n521_), .B2(new_n528_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT115), .B(new_n778_), .C1(new_n517_), .C2(new_n528_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT72), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n520_), .B(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n528_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n535_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n535_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n535_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n536_), .B1(new_n796_), .B2(KEYINPUT116), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n713_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n537_), .A2(new_n538_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n565_), .A2(new_n562_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n569_), .B(new_n800_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n570_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n605_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n794_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n537_), .B(new_n802_), .C1(new_n807_), .C2(new_n796_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT58), .B1(new_n809_), .B2(KEYINPUT117), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(new_n664_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n623_), .B1(new_n806_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n540_), .A2(new_n575_), .A3(new_n541_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n624_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n816_), .A2(new_n624_), .A3(KEYINPUT54), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n776_), .B(new_n777_), .C1(new_n815_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n713_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n355_), .B1(new_n713_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n798_), .A2(new_n803_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n716_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n805_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n804_), .A2(KEYINPUT57), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n814_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n633_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n821_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n366_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT59), .B1(new_n835_), .B2(new_n777_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n821_), .B1(new_n832_), .B2(new_n633_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  INV_X1    g637(.A(new_n777_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n366_), .A4(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n827_), .B1(new_n836_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n822_), .A2(new_n838_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n835_), .A2(KEYINPUT59), .A3(new_n777_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(KEYINPUT118), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n826_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n825_), .A2(new_n355_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n824_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  XNOR2_X1  g646(.A(KEYINPUT120), .B(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n712_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n823_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n712_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n848_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n823_), .B2(new_n623_), .ZN(new_n853_));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n855_), .B2(new_n623_), .ZN(G1342gat));
  AOI21_X1  g655(.A(G134gat), .B1(new_n823_), .B2(new_n605_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n841_), .A2(new_n844_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT121), .B(G134gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n672_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n858_), .B2(new_n860_), .ZN(G1343gat));
  NAND2_X1  g660(.A1(new_n833_), .A2(new_n834_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n364_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n777_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n575_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n215_), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n712_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n216_), .ZN(G1345gat));
  XNOR2_X1  g667(.A(KEYINPUT122), .B(KEYINPUT124), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n202_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n864_), .B2(new_n633_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n864_), .A2(new_n633_), .A3(new_n872_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n870_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n875_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n869_), .A3(new_n873_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1346gat));
  INV_X1    g678(.A(new_n864_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G162gat), .B1(new_n880_), .B2(new_n605_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n203_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(new_n882_), .ZN(G1347gat));
  NAND2_X1  g682(.A1(new_n862_), .A2(new_n776_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n437_), .A2(new_n626_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n713_), .A2(new_n330_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT125), .Z(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n713_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(G169gat), .ZN(new_n893_));
  AOI211_X1 g692(.A(KEYINPUT62), .B(new_n320_), .C1(new_n887_), .C2(new_n713_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n890_), .B1(new_n893_), .B2(new_n894_), .ZN(G1348gat));
  XNOR2_X1  g694(.A(KEYINPUT126), .B(G176gat), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n321_), .A2(KEYINPUT126), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n887_), .A2(new_n542_), .ZN(new_n898_));
  MUX2_X1   g697(.A(new_n896_), .B(new_n897_), .S(new_n898_), .Z(G1349gat));
  NAND2_X1  g698(.A1(new_n887_), .A2(new_n623_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n316_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n311_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n887_), .A2(new_n406_), .A3(new_n605_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n884_), .A2(new_n672_), .A3(new_n886_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n306_), .ZN(G1351gat));
  NAND3_X1  g704(.A1(new_n862_), .A2(new_n863_), .A3(new_n885_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n575_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n259_), .ZN(G1352gat));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n712_), .ZN(new_n909_));
  MUX2_X1   g708(.A(G204gat), .B(new_n270_), .S(new_n909_), .Z(G1353gat));
  XOR2_X1   g709(.A(KEYINPUT63), .B(G211gat), .Z(new_n911_));
  OR3_X1    g710(.A1(new_n906_), .A2(new_n633_), .A3(new_n911_), .ZN(new_n912_));
  OAI22_X1  g711(.A1(new_n906_), .A2(new_n633_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT127), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n916_), .A3(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1354gat));
  INV_X1    g717(.A(new_n906_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G218gat), .B1(new_n919_), .B2(new_n605_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n906_), .A2(new_n672_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(G218gat), .B2(new_n921_), .ZN(G1355gat));
endmodule


