//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT70), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(G1gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n211_), .B(new_n212_), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n206_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n205_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n204_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n214_), .B(new_n215_), .C1(new_n222_), .C2(new_n213_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n213_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n214_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n215_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT77), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229_));
  AOI211_X1 g028(.A(new_n229_), .B(new_n215_), .C1(new_n214_), .C2(new_n225_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n223_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G113gat), .B(G141gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(G169gat), .B(G197gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n231_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT107), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(G183gat), .A3(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT81), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n240_), .A2(new_n237_), .A3(G183gat), .A4(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT23), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n242_), .B2(KEYINPUT23), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n239_), .B(new_n241_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n246_));
  OR3_X1    g045(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n247_));
  INV_X1    g046(.A(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n246_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT78), .B(G183gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT25), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT79), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(new_n257_), .A3(KEYINPUT25), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  INV_X1    g058(.A(G183gat), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(KEYINPUT25), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .A4(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n242_), .A2(new_n265_), .A3(KEYINPUT23), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n242_), .A2(KEYINPUT23), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n238_), .A3(KEYINPUT82), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G169gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n253_), .A2(new_n262_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT84), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n272_), .B(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G127gat), .B(G134gat), .Z(new_n276_));
  XOR2_X1   g075(.A(G113gat), .B(G120gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n275_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n279_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G225gat), .A2(G233gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT3), .B1(new_n293_), .B2(KEYINPUT87), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n294_), .A2(new_n297_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n293_), .A2(new_n308_), .A3(new_n298_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n303_), .A2(new_n312_), .A3(new_n304_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n310_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n307_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n278_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n278_), .B(new_n307_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT101), .A3(new_n319_), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n316_), .A2(new_n317_), .A3(KEYINPUT101), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n290_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(KEYINPUT4), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n322_), .B1(new_n326_), .B2(new_n290_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G1gat), .B(G29gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G85gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT0), .B(G57gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT103), .ZN(new_n333_));
  INV_X1    g132(.A(new_n331_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n289_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n322_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT103), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n327_), .A2(new_n337_), .A3(new_n331_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT88), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G197gat), .B(G204gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT21), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G218gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G211gat), .ZN(new_n348_));
  INV_X1    g147(.A(G211gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G218gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G197gat), .A2(G204gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n345_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT89), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n346_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n348_), .A2(new_n350_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT90), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n357_), .A2(KEYINPUT89), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n344_), .A2(new_n345_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(KEYINPUT91), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT91), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n354_), .A2(new_n346_), .A3(new_n358_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n365_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n367_), .B(new_n371_), .C1(new_n340_), .C2(KEYINPUT88), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(new_n370_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n340_), .A2(new_n373_), .ZN(new_n374_));
  OAI22_X1  g173(.A1(new_n343_), .A2(new_n372_), .B1(new_n342_), .B2(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT92), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT28), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(KEYINPUT92), .ZN(new_n381_));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n376_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n376_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n384_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n339_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n359_), .A2(KEYINPUT91), .A3(new_n366_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT91), .B1(new_n359_), .B2(new_n366_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n272_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n260_), .A2(new_n263_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n246_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT96), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n246_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n248_), .A2(KEYINPUT22), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n248_), .A2(KEYINPUT22), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT95), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT22), .B(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n250_), .B1(new_n410_), .B2(new_n249_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n401_), .A2(new_n403_), .A3(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n250_), .A2(new_n251_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT25), .B(G183gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n259_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n268_), .A2(new_n266_), .A3(new_n247_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n416_), .A2(KEYINPUT94), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(KEYINPUT94), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n415_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n373_), .B1(new_n412_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n398_), .B(KEYINPUT20), .C1(new_n420_), .C2(new_n421_), .ZN(new_n422_));
  AOI211_X1 g221(.A(KEYINPUT97), .B(new_n373_), .C1(new_n419_), .C2(new_n412_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n395_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT98), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n371_), .A2(new_n367_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(new_n272_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n412_), .A2(new_n419_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n373_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n428_), .A2(new_n430_), .A3(KEYINPUT20), .A4(new_n394_), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT98), .B(new_n395_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G8gat), .B(G36gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  NAND4_X1  g236(.A1(new_n426_), .A2(new_n431_), .A3(new_n432_), .A4(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n428_), .A2(new_n430_), .A3(KEYINPUT20), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n395_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT97), .B1(new_n429_), .B2(new_n373_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n420_), .A2(new_n421_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n427_), .B2(new_n272_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n440_), .B1(new_n395_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n437_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n446_), .A2(KEYINPUT105), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT105), .B1(new_n446_), .B2(new_n447_), .ZN(new_n449_));
  OAI211_X1 g248(.A(KEYINPUT27), .B(new_n438_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n432_), .A2(new_n431_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT98), .B1(new_n445_), .B2(new_n395_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n447_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n438_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT27), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n454_), .A2(KEYINPUT106), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT106), .B1(new_n454_), .B2(new_n455_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n391_), .B(new_n450_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n387_), .A2(new_n390_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(KEYINPUT100), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT100), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(new_n461_), .A3(new_n438_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n326_), .A2(new_n289_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n320_), .A2(new_n321_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n331_), .B1(new_n464_), .B2(new_n290_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n335_), .A2(new_n334_), .A3(new_n322_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(KEYINPUT33), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT102), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(new_n332_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(KEYINPUT102), .A3(KEYINPUT33), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n460_), .A2(new_n462_), .A3(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n437_), .A2(KEYINPUT32), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n451_), .A2(new_n452_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n446_), .A2(new_n475_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n339_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n459_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT104), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n458_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AOI211_X1 g281(.A(KEYINPUT104), .B(new_n459_), .C1(new_n474_), .C2(new_n479_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n236_), .B(new_n288_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n456_), .A2(new_n457_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n485_), .A2(new_n450_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n459_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n288_), .A2(new_n339_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n288_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT107), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n235_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G85gat), .B(G92gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT10), .B(G99gat), .Z(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n495_), .A2(KEYINPUT9), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT6), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(G99gat), .A3(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT9), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G85gat), .A3(G92gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(new_n499_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT10), .B(G99gat), .ZN(new_n510_));
  OAI22_X1  g309(.A1(new_n505_), .A2(new_n494_), .B1(new_n510_), .B2(G106gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT65), .B1(new_n511_), .B2(new_n507_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT66), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n504_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT7), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT66), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n514_), .B1(new_n520_), .B2(new_n495_), .ZN(new_n521_));
  AOI211_X1 g320(.A(KEYINPUT8), .B(new_n494_), .C1(new_n518_), .C2(new_n504_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n513_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT67), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT67), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n513_), .B(new_n525_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n206_), .A3(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n532_), .B(KEYINPUT73), .Z(new_n533_));
  AND2_X1   g332(.A1(new_n527_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT72), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n217_), .A2(new_n221_), .A3(new_n523_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n527_), .A2(new_n536_), .A3(new_n533_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n530_), .A2(new_n531_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n534_), .B(new_n536_), .C1(KEYINPUT72), .C2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT36), .Z(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n545_), .A2(KEYINPUT36), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(new_n548_), .A3(new_n541_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n552_), .A3(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n213_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n559_));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n560_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT68), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n557_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G127gat), .B(G155gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(G183gat), .B(G211gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n566_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n557_), .B(new_n564_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n571_), .B(KEYINPUT17), .Z(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT76), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n555_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT64), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n524_), .A2(new_n564_), .A3(new_n526_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n564_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n565_), .A2(KEYINPUT12), .A3(new_n523_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n585_), .B(new_n589_), .C1(new_n587_), .C2(KEYINPUT12), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n590_), .B2(new_n584_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n588_), .B(new_n597_), .C1(new_n590_), .C2(new_n584_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n596_), .A2(KEYINPUT13), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT13), .B1(new_n596_), .B2(new_n598_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n581_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n339_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(G1gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n493_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n550_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n602_), .A2(new_n235_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n578_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT109), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n339_), .A3(new_n611_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n202_), .A2(new_n606_), .B1(new_n612_), .B2(G1gat), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n606_), .A2(new_n202_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT108), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n606_), .A2(KEYINPUT108), .A3(new_n202_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT110), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(G1324gat));
  INV_X1    g419(.A(new_n486_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n608_), .A2(new_n621_), .A3(new_n611_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n493_), .A2(new_n603_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n209_), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n625_), .A2(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(G1325gat));
  NAND2_X1  g430(.A1(new_n608_), .A2(new_n611_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G15gat), .B1(new_n632_), .B2(new_n288_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT41), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n627_), .A2(G15gat), .A3(new_n288_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1326gat));
  OAI21_X1  g435(.A(G22gat), .B1(new_n632_), .B2(new_n487_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT42), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n487_), .A2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n627_), .B2(new_n639_), .ZN(G1327gat));
  XOR2_X1   g439(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n641_));
  XOR2_X1   g440(.A(new_n554_), .B(KEYINPUT111), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n484_), .A2(new_n489_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n338_), .A2(new_n336_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n467_), .A2(new_n337_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n478_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n476_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n332_), .A2(new_n470_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n467_), .A2(KEYINPUT102), .A3(KEYINPUT33), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n467_), .B2(KEYINPUT33), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n461_), .B1(new_n453_), .B2(new_n438_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n647_), .B1(new_n653_), .B2(new_n462_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT104), .B1(new_n654_), .B2(new_n459_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n480_), .A2(new_n481_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n458_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n236_), .B1(new_n657_), .B2(new_n288_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n642_), .B1(new_n643_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n492_), .A2(new_n489_), .A3(new_n484_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n554_), .A2(KEYINPUT43), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n659_), .A2(KEYINPUT43), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n609_), .A2(new_n579_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n641_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n663_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n660_), .B2(new_n642_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n661_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n665_), .C1(new_n667_), .C2(new_n669_), .ZN(new_n670_));
  AND4_X1   g469(.A1(G29gat), .A2(new_n664_), .A3(new_n339_), .A4(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n602_), .A2(new_n578_), .A3(new_n550_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n493_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n339_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n671_), .A2(new_n675_), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n664_), .A2(new_n621_), .A3(new_n670_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n486_), .A2(G36gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n673_), .A2(KEYINPUT45), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT45), .B1(new_n673_), .B2(new_n680_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n678_), .B(new_n683_), .C1(KEYINPUT113), .C2(KEYINPUT46), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1329gat));
  NAND4_X1  g487(.A1(new_n664_), .A2(G43gat), .A3(new_n287_), .A4(new_n670_), .ZN(new_n689_));
  INV_X1    g488(.A(G43gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n673_), .B2(new_n288_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g492(.A1(G50gat), .A2(new_n664_), .A3(new_n459_), .A4(new_n670_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G50gat), .B1(new_n674_), .B2(new_n459_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1331gat));
  NAND2_X1  g495(.A1(new_n602_), .A2(new_n235_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n579_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n608_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G57gat), .B1(new_n699_), .B2(new_n604_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n235_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n580_), .A3(new_n602_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n604_), .A2(G57gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1332gat));
  OAI21_X1  g504(.A(G64gat), .B1(new_n699_), .B2(new_n486_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT48), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n486_), .A2(G64gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n703_), .B2(new_n708_), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n699_), .B2(new_n288_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT49), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n288_), .A2(G71gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n703_), .B2(new_n712_), .ZN(G1334gat));
  OAI21_X1  g512(.A(G78gat), .B1(new_n699_), .B2(new_n487_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT50), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n487_), .A2(G78gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n703_), .B2(new_n716_), .ZN(G1335gat));
  NOR3_X1   g516(.A1(new_n662_), .A2(new_n578_), .A3(new_n697_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n718_), .A2(KEYINPUT114), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(KEYINPUT114), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n339_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G85gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n601_), .A2(new_n578_), .A3(new_n550_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n702_), .A2(new_n723_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n724_), .A2(G85gat), .A3(new_n604_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1336gat));
  NAND3_X1  g525(.A1(new_n719_), .A2(new_n621_), .A3(new_n720_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G92gat), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n724_), .A2(G92gat), .A3(new_n486_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1337gat));
  NAND2_X1  g529(.A1(new_n718_), .A2(new_n287_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G99gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n724_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n287_), .A3(new_n496_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT51), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n497_), .A3(new_n459_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n697_), .A2(new_n578_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n459_), .B(new_n741_), .C1(new_n667_), .C2(new_n669_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(G106gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G106gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n740_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n740_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  OAI211_X1 g549(.A(new_n223_), .B(new_n234_), .C1(new_n228_), .C2(new_n230_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n214_), .B(new_n227_), .C1(new_n222_), .C2(new_n213_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n234_), .B1(new_n226_), .B2(new_n215_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n598_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT119), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n598_), .A2(new_n755_), .A3(KEYINPUT119), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n590_), .B2(new_n584_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n590_), .A2(new_n584_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n585_), .A2(new_n589_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n564_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n521_), .A2(new_n522_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n525_), .B1(new_n767_), .B2(new_n513_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n526_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT12), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n765_), .A2(new_n772_), .A3(KEYINPUT55), .A4(new_n583_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n763_), .A2(new_n764_), .A3(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n595_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n595_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n760_), .B(new_n761_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n774_), .A2(new_n595_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n775_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n761_), .B1(new_n783_), .B2(new_n760_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n555_), .B1(new_n779_), .B2(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n701_), .A2(new_n598_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n788_));
  NAND3_X1  g587(.A1(new_n780_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n775_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n780_), .B2(new_n788_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n786_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n596_), .A2(new_n598_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n755_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n607_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT121), .B(new_n785_), .C1(new_n795_), .C2(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT57), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n780_), .A2(new_n788_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT117), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n775_), .A3(new_n789_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n802_), .A2(new_n786_), .B1(new_n793_), .B2(new_n755_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n803_), .B2(new_n607_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT121), .B1(new_n804_), .B2(new_n785_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n579_), .B1(new_n798_), .B2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n554_), .A2(new_n235_), .A3(new_n578_), .A4(new_n601_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(KEYINPUT54), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n806_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n486_), .A2(new_n287_), .A3(new_n487_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n816_), .A2(KEYINPUT59), .A3(new_n604_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n813_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT118), .B(new_n799_), .C1(new_n803_), .C2(new_n607_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n785_), .A4(new_n797_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n823_), .B2(new_n579_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n824_), .A2(new_n604_), .A3(new_n816_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n818_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n815_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT123), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OR3_X1    g628(.A1(new_n824_), .A2(new_n604_), .A3(new_n816_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT59), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n814_), .A2(new_n817_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT122), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n831_), .A2(new_n832_), .A3(new_n834_), .A4(new_n818_), .ZN(new_n835_));
  INV_X1    g634(.A(G113gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n235_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n829_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n830_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n825_), .A2(KEYINPUT120), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n701_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n836_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n838_), .A2(new_n843_), .ZN(G1340gat));
  NAND3_X1  g643(.A1(new_n831_), .A2(new_n834_), .A3(new_n818_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G120gat), .B1(new_n845_), .B2(new_n601_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n840_), .A2(new_n841_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848_));
  AOI21_X1  g647(.A(G120gat), .B1(new_n602_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n848_), .B2(G120gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT124), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  AND4_X1   g650(.A1(KEYINPUT124), .A2(new_n840_), .A3(new_n841_), .A4(new_n850_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n846_), .B1(new_n851_), .B2(new_n852_), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n579_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n829_), .A2(new_n835_), .A3(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n840_), .A2(new_n578_), .A3(new_n841_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n854_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n554_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n829_), .A2(new_n835_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n840_), .A2(new_n607_), .A3(new_n841_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n860_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1343gat));
  NAND3_X1  g664(.A1(new_n486_), .A2(new_n288_), .A3(new_n459_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n824_), .A2(new_n604_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n701_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n602_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n578_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n872_), .A2(KEYINPUT125), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(KEYINPUT125), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n867_), .B2(new_n607_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n642_), .A2(G162gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n867_), .B2(new_n880_), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n621_), .A2(new_n488_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n459_), .B(new_n882_), .C1(new_n806_), .C2(new_n813_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n248_), .B1(new_n883_), .B2(new_n701_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n701_), .A2(new_n410_), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT126), .Z(new_n888_));
  NAND2_X1  g687(.A1(new_n883_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(G1348gat));
  OR2_X1    g689(.A1(new_n824_), .A2(new_n459_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n891_), .A2(new_n249_), .A3(new_n601_), .A4(new_n882_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G176gat), .B1(new_n883_), .B2(new_n602_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1349gat));
  OR3_X1    g693(.A1(new_n891_), .A2(new_n579_), .A3(new_n882_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n579_), .A2(new_n414_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n895_), .A2(new_n254_), .B1(new_n883_), .B2(new_n896_), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n883_), .A2(new_n259_), .A3(new_n607_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n883_), .A2(new_n555_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n263_), .ZN(G1351gat));
  NAND3_X1  g699(.A1(new_n621_), .A2(new_n288_), .A3(new_n391_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n824_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n701_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n602_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g705(.A1(new_n902_), .A2(new_n578_), .ZN(new_n907_));
  AND2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT127), .B1(new_n907_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n907_), .A2(new_n909_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n907_), .A2(KEYINPUT127), .A3(new_n910_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1354gat));
  NAND3_X1  g714(.A1(new_n902_), .A2(new_n347_), .A3(new_n607_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n824_), .A2(new_n554_), .A3(new_n901_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n347_), .ZN(G1355gat));
endmodule


