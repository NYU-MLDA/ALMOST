//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G169gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT90), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n206_), .B2(new_n203_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n207_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT24), .B1(new_n202_), .B2(new_n203_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n222_), .B1(new_n223_), .B2(new_n220_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n208_), .A2(new_n211_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n216_), .A2(KEYINPUT26), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .A4(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n219_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G204gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G197gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G204gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n236_), .A2(new_n237_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT21), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G211gat), .B(G218gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n240_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(KEYINPUT21), .A3(new_n245_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n234_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT20), .ZN(new_n253_));
  INV_X1    g052(.A(new_n251_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n255_), .A2(new_n215_), .A3(KEYINPUT25), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n255_), .B2(new_n228_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT82), .B(G190gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n230_), .B1(new_n258_), .B2(new_n229_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n224_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n258_), .A2(G183gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n226_), .A2(new_n262_), .A3(new_n227_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n204_), .B1(new_n205_), .B2(new_n203_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n260_), .A2(new_n261_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n253_), .B1(new_n254_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n252_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT94), .ZN(new_n271_));
  INV_X1    g070(.A(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n251_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n254_), .A2(new_n219_), .A3(new_n233_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT20), .ZN(new_n275_));
  INV_X1    g074(.A(new_n269_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT94), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n252_), .A2(new_n266_), .A3(new_n278_), .A4(new_n269_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n271_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT18), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT32), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n252_), .A2(new_n266_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n276_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT91), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n269_), .B1(new_n252_), .B2(new_n266_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT91), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT20), .A4(new_n269_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .A4(new_n285_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n300_), .A2(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT86), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n299_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n300_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n302_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n298_), .A2(KEYINPUT1), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n298_), .B1(new_n296_), .B2(KEYINPUT1), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(KEYINPUT85), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT85), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n315_), .B(new_n298_), .C1(new_n296_), .C2(KEYINPUT1), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n311_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n309_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n323_));
  INV_X1    g122(.A(new_n319_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G113gat), .B(G120gat), .Z(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n309_), .B2(new_n317_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT92), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(new_n328_), .B2(KEYINPUT4), .ZN(new_n334_));
  INV_X1    g133(.A(new_n318_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n335_), .A2(KEYINPUT93), .A3(new_n336_), .A4(new_n327_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n322_), .A2(new_n328_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n334_), .B(new_n337_), .C1(new_n338_), .C2(new_n336_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n332_), .B1(new_n339_), .B2(new_n331_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT0), .B(G57gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  AOI211_X1 g145(.A(new_n344_), .B(new_n332_), .C1(new_n339_), .C2(new_n331_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n287_), .B(new_n295_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n339_), .A2(new_n331_), .ZN(new_n349_));
  OAI211_X1 g148(.A(KEYINPUT33), .B(new_n344_), .C1(new_n349_), .C2(new_n332_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n284_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n294_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n355_));
  AOI211_X1 g154(.A(KEYINPUT91), .B(new_n269_), .C1(new_n252_), .C2(new_n266_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n290_), .A2(new_n284_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n344_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n339_), .B2(new_n331_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n348_), .B1(new_n353_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n318_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n364_), .B(KEYINPUT28), .Z(new_n365_));
  OAI21_X1  g164(.A(new_n251_), .B1(new_n318_), .B2(new_n363_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n366_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(G78gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G106gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G22gat), .B(G50gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n367_), .A2(new_n368_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n358_), .A2(KEYINPUT27), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n280_), .A2(new_n354_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n280_), .A2(KEYINPUT97), .A3(new_n354_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT27), .B1(new_n357_), .B2(new_n358_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT96), .ZN(new_n390_));
  OR3_X1    g189(.A1(new_n346_), .A2(new_n347_), .A3(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n378_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n362_), .A2(KEYINPUT95), .A3(new_n378_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n381_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397_));
  INV_X1    g196(.A(G43gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n265_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(new_n327_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(G15gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT30), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT31), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n401_), .B(new_n406_), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n378_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n410_));
  INV_X1    g209(.A(new_n388_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n385_), .A2(new_n386_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n410_), .B(new_n411_), .C1(new_n412_), .C2(new_n382_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT98), .B1(new_n387_), .B2(new_n388_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n409_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n391_), .A2(new_n392_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(new_n408_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n396_), .A2(new_n408_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G113gat), .B(G141gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT80), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G169gat), .B(G197gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G229gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G29gat), .B(G36gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G43gat), .B(G50gat), .Z(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G43gat), .B(G50gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT77), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(KEYINPUT77), .A3(new_n431_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G1gat), .B(G8gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT73), .ZN(new_n437_));
  INV_X1    g236(.A(G1gat), .ZN(new_n438_));
  OR2_X1    g237(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT14), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n437_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n440_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(G1gat), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(KEYINPUT73), .A3(KEYINPUT14), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G15gat), .B(G22gat), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n436_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n436_), .ZN(new_n452_));
  AOI211_X1 g251(.A(new_n449_), .B(new_n452_), .C1(new_n443_), .C2(new_n447_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n435_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n441_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT73), .B1(new_n446_), .B2(KEYINPUT14), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n450_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n452_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n448_), .A2(new_n450_), .A3(new_n436_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(KEYINPUT78), .A3(new_n435_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n456_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n462_), .B2(new_n435_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n429_), .A2(KEYINPUT77), .A3(new_n431_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(new_n432_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n460_), .A2(new_n468_), .A3(KEYINPUT79), .A4(new_n461_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n425_), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n425_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n429_), .A2(new_n431_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT15), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n429_), .A2(KEYINPUT15), .A3(new_n431_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n477_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n478_));
  AOI211_X1 g277(.A(new_n472_), .B(new_n478_), .C1(new_n456_), .C2(new_n463_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n424_), .B1(new_n471_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n478_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n464_), .A2(new_n425_), .A3(new_n481_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n456_), .A2(new_n463_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n482_), .B(new_n423_), .C1(new_n483_), .C2(new_n425_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n419_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G85gat), .ZN(new_n488_));
  INV_X1    g287(.A(G92gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT65), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n490_), .A2(KEYINPUT9), .B1(new_n488_), .B2(new_n489_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT9), .ZN(new_n492_));
  OAI211_X1 g291(.A(KEYINPUT65), .B(new_n492_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n494_), .B(new_n500_), .C1(new_n506_), .C2(G106gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(G85gat), .B(G92gat), .Z(new_n508_));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509_));
  INV_X1    g308(.A(G99gat), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n372_), .A4(KEYINPUT66), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n512_));
  OAI22_X1  g311(.A1(new_n512_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(KEYINPUT67), .B(new_n508_), .C1(new_n514_), .C2(new_n499_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(KEYINPUT68), .A3(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n515_), .A2(KEYINPUT68), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT68), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n519_), .B(new_n508_), .C1(new_n514_), .C2(new_n499_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT8), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n507_), .B(new_n517_), .C1(new_n518_), .C2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G78gat), .Z(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT12), .B1(new_n522_), .B2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n522_), .A2(new_n529_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n521_), .B1(KEYINPUT68), .B2(new_n515_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n507_), .A2(new_n517_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n515_), .A2(KEYINPUT68), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(KEYINPUT8), .A3(new_n520_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n539_), .A2(KEYINPUT69), .A3(new_n507_), .A4(new_n517_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n529_), .A2(KEYINPUT12), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n532_), .A2(new_n533_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n533_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n529_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n507_), .A2(new_n517_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n547_), .B2(new_n539_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n545_), .B1(new_n548_), .B2(new_n531_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT5), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n544_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT13), .Z(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n462_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n546_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n562_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n562_), .A2(KEYINPUT75), .A3(new_n569_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT76), .ZN(new_n577_));
  INV_X1    g376(.A(new_n477_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n537_), .A2(new_n578_), .A3(new_n540_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n583_));
  INV_X1    g382(.A(new_n522_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n584_), .B2(new_n473_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT71), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n579_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n585_), .B2(new_n579_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n598_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n577_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n487_), .A2(new_n559_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT99), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(KEYINPUT99), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n438_), .A3(new_n417_), .A4(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n597_), .A2(new_n612_), .A3(new_n599_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n419_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n559_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n576_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n486_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n416_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n609_), .A2(new_n610_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n621_), .A3(new_n622_), .ZN(G1324gat));
  AND2_X1   g422(.A1(new_n413_), .A2(new_n414_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n625_), .A2(new_n445_), .A3(new_n444_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n607_), .A2(new_n608_), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G8gat), .B1(new_n620_), .B2(new_n625_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(KEYINPUT101), .A2(KEYINPUT39), .ZN(new_n629_));
  AND2_X1   g428(.A1(KEYINPUT101), .A2(KEYINPUT39), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n629_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n627_), .A2(new_n631_), .A3(KEYINPUT40), .A4(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  OAI21_X1  g436(.A(G15gat), .B1(new_n620_), .B2(new_n408_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT102), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n640_), .B(G15gat), .C1(new_n620_), .C2(new_n408_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n639_), .A2(KEYINPUT41), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n606_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT41), .B1(new_n639_), .B2(new_n641_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT103), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n645_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(new_n642_), .A3(new_n648_), .A4(new_n643_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n620_), .B2(new_n378_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n378_), .A2(G22gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n605_), .B2(new_n653_), .ZN(G1327gat));
  NAND3_X1  g453(.A1(new_n577_), .A2(new_n485_), .A3(new_n559_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n602_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n600_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT43), .B1(new_n419_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n380_), .A2(new_n379_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n407_), .B1(new_n660_), .B2(new_n395_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n415_), .A2(new_n418_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n659_), .B(new_n603_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n655_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT44), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n417_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G29gat), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  INV_X1    g468(.A(new_n577_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n615_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n669_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n577_), .A2(KEYINPUT104), .A3(new_n615_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n617_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n487_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n416_), .A2(G29gat), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT105), .Z(new_n677_));
  OAI21_X1  g476(.A(new_n668_), .B1(new_n675_), .B2(new_n677_), .ZN(G1328gat));
  NOR2_X1   g477(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT107), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n624_), .B1(new_n664_), .B2(KEYINPUT44), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n682_), .B(new_n655_), .C1(new_n658_), .C2(new_n663_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G36gat), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n675_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n625_), .A2(G36gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT45), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  AND4_X1   g486(.A1(KEYINPUT45), .A2(new_n487_), .A3(new_n674_), .A4(new_n686_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n684_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n680_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n691_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n680_), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n693_), .B(new_n694_), .C1(new_n684_), .C2(new_n689_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1329gat));
  OAI21_X1  g495(.A(new_n398_), .B1(new_n675_), .B2(new_n408_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n665_), .A2(G43gat), .A3(new_n407_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n683_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT47), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n699_), .B(new_n703_), .C1(new_n700_), .C2(new_n683_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1330gat));
  INV_X1    g504(.A(G50gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n665_), .A2(new_n409_), .A3(new_n666_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(KEYINPUT109), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(KEYINPUT109), .B2(new_n707_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n685_), .A2(new_n706_), .A3(new_n409_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1331gat));
  NOR2_X1   g510(.A1(new_n419_), .A2(new_n485_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n712_), .A2(new_n617_), .A3(new_n604_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n417_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n616_), .A2(new_n486_), .A3(new_n617_), .A4(new_n670_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n416_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1332gat));
  OAI21_X1  g517(.A(G64gat), .B1(new_n716_), .B2(new_n625_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT48), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n625_), .A2(G64gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT110), .Z(new_n722_));
  NAND2_X1  g521(.A1(new_n713_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n716_), .B2(new_n408_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT49), .ZN(new_n726_));
  INV_X1    g525(.A(G71gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n713_), .A2(new_n727_), .A3(new_n407_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1334gat));
  OAI21_X1  g528(.A(G78gat), .B1(new_n716_), .B2(new_n378_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT50), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n713_), .A2(new_n370_), .A3(new_n409_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1335gat));
  NAND3_X1  g532(.A1(new_n577_), .A2(new_n617_), .A3(new_n486_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n416_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n559_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n712_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n488_), .A3(new_n417_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1336gat));
  AOI21_X1  g540(.A(G92gat), .B1(new_n739_), .B2(new_n624_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n624_), .A2(G92gat), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT111), .Z(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n735_), .B2(new_n744_), .ZN(G1337gat));
  NOR2_X1   g544(.A1(new_n408_), .A2(new_n506_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT112), .B1(new_n739_), .B2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n736_), .A2(new_n408_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n510_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n372_), .A3(new_n409_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n735_), .A2(new_n409_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G106gat), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT52), .B(new_n372_), .C1(new_n735_), .C2(new_n409_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n464_), .A2(new_n472_), .A3(new_n481_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n424_), .C1(new_n483_), .C2(new_n472_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n484_), .A2(new_n761_), .A3(new_n555_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n533_), .B1(new_n532_), .B2(new_n543_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n544_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n532_), .A2(KEYINPUT55), .A3(new_n533_), .A4(new_n543_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n554_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n762_), .B1(new_n767_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n547_), .A2(new_n546_), .A3(new_n539_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n522_), .A2(new_n529_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT12), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AND4_X1   g575(.A1(new_n533_), .A2(new_n543_), .A3(new_n773_), .A4(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n543_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n548_), .B2(KEYINPUT12), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n545_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n777_), .B1(KEYINPUT55), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n766_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n553_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n769_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT58), .B1(new_n772_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n759_), .B1(new_n785_), .B2(new_n657_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n553_), .B(new_n771_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n762_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n767_), .A2(new_n768_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT115), .A3(new_n603_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n772_), .A2(new_n784_), .A3(KEYINPUT58), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n786_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n484_), .A2(new_n761_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n558_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n485_), .A2(new_n555_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(KEYINPUT56), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n767_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n767_), .A2(new_n801_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n798_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n796_), .B1(new_n805_), .B2(new_n615_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n798_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n767_), .A2(new_n801_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n485_), .A3(new_n555_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n809_), .B2(new_n803_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT57), .A3(new_n671_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n758_), .B1(new_n795_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n786_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(KEYINPUT116), .A3(new_n806_), .A4(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n618_), .A3(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n670_), .A2(new_n486_), .A3(new_n559_), .A4(new_n657_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT54), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n415_), .A2(new_n417_), .A3(new_n407_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(G113gat), .B1(new_n822_), .B2(new_n485_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n577_), .B1(new_n795_), .B2(new_n812_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n818_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n820_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n485_), .A2(G113gat), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT117), .Z(new_n832_));
  AOI21_X1  g631(.A(new_n823_), .B1(new_n830_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n834_));
  AOI21_X1  g633(.A(G120gat), .B1(new_n617_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n834_), .B2(G120gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n822_), .A2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT118), .ZN(new_n838_));
  OAI21_X1  g637(.A(G120gat), .B1(new_n829_), .B2(new_n559_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n821_), .B2(new_n577_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n843_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n618_), .A2(new_n841_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n844_), .A2(new_n845_), .B1(new_n830_), .B2(new_n846_), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n821_), .B2(new_n671_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n850_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n657_), .A2(new_n848_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n851_), .A2(new_n852_), .B1(new_n830_), .B2(new_n853_), .ZN(G1343gat));
  NOR4_X1   g653(.A1(new_n624_), .A2(new_n378_), .A3(new_n416_), .A4(new_n407_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n819_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n485_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n617_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g660(.A1(new_n856_), .A2(new_n577_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  AOI21_X1  g663(.A(G162gat), .B1(new_n857_), .B2(new_n615_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n603_), .A2(G162gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT121), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n857_), .B2(new_n867_), .ZN(G1347gat));
  NAND2_X1  g667(.A1(new_n624_), .A2(new_n418_), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT122), .Z(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n409_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n826_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872_), .B2(new_n486_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n872_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n206_), .A3(new_n485_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n874_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n877_), .A3(new_n878_), .ZN(G1348gat));
  OAI21_X1  g678(.A(new_n203_), .B1(new_n872_), .B2(new_n559_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n880_), .A2(KEYINPUT123), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(KEYINPUT123), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n409_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n870_), .A2(new_n203_), .A3(new_n559_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n881_), .A2(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1349gat));
  INV_X1    g684(.A(new_n870_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n670_), .A3(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G183gat), .B1(new_n887_), .B2(new_n888_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n618_), .A2(new_n228_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n889_), .A2(new_n890_), .B1(new_n876_), .B2(new_n891_), .ZN(G1350gat));
  NAND4_X1  g691(.A1(new_n876_), .A2(new_n230_), .A3(new_n231_), .A4(new_n615_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n876_), .A2(new_n603_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(G190gat), .ZN(new_n896_));
  AOI211_X1 g695(.A(KEYINPUT125), .B(new_n216_), .C1(new_n876_), .C2(new_n603_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n893_), .B1(new_n896_), .B2(new_n897_), .ZN(G1351gat));
  NAND3_X1  g697(.A1(new_n624_), .A2(new_n408_), .A3(new_n393_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n485_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n617_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n576_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1354gat));
  NAND3_X1  g708(.A1(new_n900_), .A2(G218gat), .A3(new_n603_), .ZN(new_n910_));
  INV_X1    g709(.A(G218gat), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n671_), .B(new_n899_), .C1(new_n816_), .C2(new_n818_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n900_), .A2(new_n913_), .A3(new_n615_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n910_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  OAI211_X1 g717(.A(KEYINPUT127), .B(new_n910_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1355gat));
endmodule


