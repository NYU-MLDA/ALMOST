//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT24), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n208_), .B2(KEYINPUT24), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT25), .B(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT26), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT81), .B1(new_n211_), .B2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n210_), .B(new_n212_), .C1(new_n213_), .C2(KEYINPUT81), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n215_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n215_), .A2(KEYINPUT23), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n209_), .B(new_n214_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n203_), .A2(KEYINPUT22), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT83), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n204_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G169gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n225_), .B1(new_n224_), .B2(new_n229_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n223_), .B(new_n207_), .C1(new_n227_), .C2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n218_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n216_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n215_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n215_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n231_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G169gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n204_), .B(new_n226_), .C1(new_n242_), .C2(new_n225_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n223_), .B1(new_n243_), .B2(new_n207_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n222_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n222_), .B(KEYINPUT85), .C1(new_n241_), .C2(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G71gat), .B(G99gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G43gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n249_), .B(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G127gat), .B(G134gat), .Z(new_n253_));
  XOR2_X1   g052(.A(G113gat), .B(G120gat), .Z(new_n254_));
  XOR2_X1   g053(.A(new_n253_), .B(new_n254_), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n252_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(G15gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT30), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT31), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n256_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G228gat), .A2(G233gat), .ZN(new_n264_));
  INV_X1    g063(.A(G78gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G106gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G22gat), .B(G50gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT87), .Z(new_n273_));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT1), .Z(new_n275_));
  AND2_X1   g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT86), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G141gat), .A2(G148gat), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n276_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(G141gat), .ZN(new_n286_));
  INV_X1    g085(.A(G148gat), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT3), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT3), .B1(new_n286_), .B2(new_n287_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n285_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n278_), .A2(new_n280_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT88), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n278_), .A2(new_n280_), .A3(KEYINPUT88), .A4(new_n291_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n290_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT89), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n273_), .A2(new_n274_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT90), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT89), .ZN(new_n300_));
  AOI211_X1 g099(.A(new_n300_), .B(new_n290_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n294_), .A2(new_n295_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n290_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT89), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT90), .B(new_n298_), .C1(new_n301_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n284_), .B1(new_n299_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT28), .B1(new_n307_), .B2(KEYINPUT29), .ZN(new_n308_));
  XOR2_X1   g107(.A(G211gat), .B(G218gat), .Z(new_n309_));
  INV_X1    g108(.A(G204gat), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n310_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(G197gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT92), .B1(new_n310_), .B2(G197gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n309_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT91), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n310_), .B2(G197gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n312_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n318_), .A2(new_n310_), .A3(G197gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT21), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n314_), .A2(KEYINPUT93), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(KEYINPUT93), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT21), .A4(new_n309_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n298_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n283_), .B1(new_n330_), .B2(new_n305_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n327_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n308_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n308_), .B2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n271_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n336_), .A3(new_n270_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n255_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n330_), .A2(new_n305_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n284_), .ZN(new_n351_));
  AOI211_X1 g150(.A(new_n255_), .B(new_n283_), .C1(new_n330_), .C2(new_n305_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n348_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n307_), .A2(new_n255_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n331_), .A2(new_n349_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT4), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n354_), .B1(new_n351_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n357_), .A3(new_n354_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n347_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G8gat), .B(G36gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT99), .ZN(new_n367_));
  XOR2_X1   g166(.A(G64gat), .B(G92gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n369_), .B(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n323_), .A2(new_n326_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n205_), .A2(new_n207_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n213_), .A2(new_n210_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n235_), .A2(new_n237_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  INV_X1    g183(.A(new_n221_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n238_), .B1(new_n219_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n207_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n242_), .B2(new_n204_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n384_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n391_), .A2(new_n386_), .A3(KEYINPUT97), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n383_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n375_), .B1(new_n393_), .B2(new_n327_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n374_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT95), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  NOR2_X1   g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n249_), .A2(new_n327_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n381_), .A2(new_n382_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n373_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n372_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT27), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT20), .B(new_n401_), .C1(new_n393_), .C2(new_n327_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n327_), .B2(new_n249_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n401_), .B1(new_n374_), .B2(new_n394_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n372_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n372_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n395_), .A2(new_n399_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n401_), .A2(KEYINPUT20), .ZN(new_n417_));
  INV_X1    g216(.A(new_n390_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n392_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n418_), .A2(new_n419_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n417_), .B1(new_n420_), .B2(new_n373_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n402_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(new_n422_), .A3(new_n413_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n415_), .A2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n407_), .A2(new_n414_), .B1(new_n424_), .B2(new_n408_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n263_), .A2(new_n343_), .A3(new_n365_), .A4(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n365_), .A2(new_n342_), .A3(new_n425_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n354_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n347_), .B1(new_n353_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n351_), .B2(new_n359_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n358_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n424_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT33), .B1(new_n355_), .B2(new_n361_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n347_), .A2(KEYINPUT33), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT100), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n439_), .A2(new_n361_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n439_), .B2(new_n361_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n361_), .A2(new_n363_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n348_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n355_), .A2(new_n361_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n372_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT103), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT103), .B(new_n449_), .C1(new_n400_), .C2(new_n406_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n449_), .B(KEYINPUT101), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n452_), .A2(new_n453_), .B1(new_n454_), .B2(new_n412_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n437_), .A2(new_n443_), .B1(new_n447_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n428_), .B1(new_n456_), .B2(new_n342_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n427_), .B1(new_n457_), .B2(new_n262_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT10), .B(G99gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT64), .B(G106gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G99gat), .A3(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G85gat), .A3(G92gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(G85gat), .B(G92gat), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n461_), .A2(new_n466_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT65), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n476_));
  INV_X1    g275(.A(new_n474_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n473_), .A2(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n466_), .A2(KEYINPUT67), .ZN(new_n479_));
  OR2_X1    g278(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(KEYINPUT65), .A3(new_n474_), .A4(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n463_), .A2(new_n465_), .A3(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n478_), .A2(new_n479_), .A3(new_n482_), .A4(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n472_), .B1(new_n485_), .B2(new_n469_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n473_), .A2(new_n475_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n477_), .A2(new_n476_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n487_), .A2(new_n482_), .A3(new_n466_), .A4(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n489_), .A2(new_n472_), .A3(new_n469_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n471_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G36gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G29gat), .ZN(new_n493_));
  INV_X1    g292(.A(G29gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G36gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT71), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n495_), .A3(KEYINPUT71), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n498_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n496_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n500_), .A2(new_n503_), .A3(KEYINPUT15), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT15), .B1(new_n500_), .B2(new_n503_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n491_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT34), .Z(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n500_), .A2(new_n503_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n513_), .B(new_n471_), .C1(new_n486_), .C2(new_n490_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n509_), .A2(new_n510_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n507_), .A2(new_n512_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(new_n514_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n511_), .ZN(new_n519_));
  AOI211_X1 g318(.A(KEYINPUT72), .B(new_n512_), .C1(new_n507_), .C2(new_n514_), .ZN(new_n520_));
  OAI211_X1 g319(.A(KEYINPUT74), .B(new_n516_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G190gat), .B(G218gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT73), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n521_), .A2(new_n522_), .A3(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n526_), .B(new_n516_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n522_), .B1(new_n521_), .B2(new_n527_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n458_), .A2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n534_), .A2(KEYINPUT104), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(KEYINPUT104), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n539_));
  XOR2_X1   g338(.A(G71gat), .B(G78gat), .Z(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n540_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n491_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n491_), .A2(new_n545_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT12), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n544_), .B(KEYINPUT68), .Z(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n547_), .B(new_n549_), .C1(new_n491_), .C2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n547_), .A2(new_n548_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(new_n554_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G120gat), .B(G148gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G176gat), .B(G204gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(KEYINPUT69), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n566_), .A2(KEYINPUT13), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(KEYINPUT13), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT75), .B(G8gat), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT14), .B1(new_n571_), .B2(new_n202_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G1gat), .B(G8gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT76), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT77), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(new_n544_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n544_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT17), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT78), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n582_), .A3(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n579_), .A2(new_n550_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n586_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n550_), .B2(new_n579_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT80), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n576_), .B2(new_n513_), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n576_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT79), .B1(new_n576_), .B2(new_n513_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n576_), .A2(new_n513_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n604_), .B2(new_n595_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n605_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n570_), .A2(new_n594_), .A3(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n537_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n202_), .B1(new_n613_), .B2(new_n447_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n458_), .A2(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n521_), .A2(new_n527_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT36), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(KEYINPUT37), .A3(new_n529_), .A4(new_n528_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n594_), .A2(new_n622_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n615_), .A2(new_n569_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n202_), .A3(new_n447_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT38), .Z(new_n626_));
  NOR2_X1   g425(.A1(new_n614_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT105), .ZN(G1324gat));
  INV_X1    g427(.A(new_n425_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(new_n629_), .A3(new_n571_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n629_), .B(new_n612_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(new_n632_), .A3(G8gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G8gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g435(.A1(new_n624_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n613_), .A2(new_n263_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT41), .B1(new_n638_), .B2(G15gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n624_), .A2(new_n642_), .A3(new_n342_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n613_), .A2(new_n342_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(G22gat), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT42), .B(new_n642_), .C1(new_n613_), .C2(new_n342_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(G1327gat));
  NAND3_X1  g447(.A1(new_n569_), .A2(new_n533_), .A3(new_n594_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n615_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n447_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n446_), .A2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n351_), .A2(new_n352_), .A3(new_n359_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n307_), .A2(new_n359_), .A3(new_n255_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n429_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n438_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n363_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT100), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n424_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n439_), .A2(new_n361_), .A3(new_n440_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n655_), .A2(new_n662_), .A3(new_n663_), .A4(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n455_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n342_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n365_), .A2(new_n342_), .A3(new_n425_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n262_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n426_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n621_), .A2(KEYINPUT43), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n617_), .A2(KEYINPUT106), .A3(new_n620_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT106), .B1(new_n617_), .B2(new_n620_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n458_), .C2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n669_), .B2(new_n426_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n673_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n569_), .A2(new_n594_), .A3(new_n610_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n365_), .A2(new_n494_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n653_), .B1(new_n687_), .B2(new_n688_), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n629_), .A3(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G36gat), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n629_), .A2(KEYINPUT108), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n629_), .A2(KEYINPUT108), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n652_), .A2(new_n492_), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT45), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1329gat));
  NAND4_X1  g498(.A1(new_n685_), .A2(G43gat), .A3(new_n263_), .A4(new_n686_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n651_), .A2(new_n262_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(G43gat), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g502(.A1(new_n685_), .A2(new_n342_), .A3(new_n686_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G50gat), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n651_), .A2(G50gat), .A3(new_n343_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT109), .ZN(G1331gat));
  INV_X1    g507(.A(G57gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n594_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n569_), .A2(new_n610_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n537_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n712_), .B2(new_n447_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n670_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n623_), .ZN(new_n715_));
  NOR4_X1   g514(.A1(new_n714_), .A2(G57gat), .A3(new_n365_), .A4(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n713_), .A2(new_n716_), .ZN(G1332gat));
  NOR2_X1   g516(.A1(new_n714_), .A2(new_n715_), .ZN(new_n718_));
  INV_X1    g517(.A(G64gat), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n694_), .A2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT110), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n712_), .A2(new_n694_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(G64gat), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT48), .B(new_n719_), .C1(new_n712_), .C2(new_n694_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n718_), .A2(new_n728_), .A3(new_n263_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n712_), .A2(new_n263_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G71gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT49), .B(new_n728_), .C1(new_n712_), .C2(new_n263_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1334gat));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n265_), .A3(new_n342_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n712_), .A2(new_n342_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G78gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT50), .B(new_n265_), .C1(new_n712_), .C2(new_n342_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1335gat));
  NOR3_X1   g539(.A1(new_n714_), .A2(new_n532_), .A3(new_n710_), .ZN(new_n741_));
  INV_X1    g540(.A(G85gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n447_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n711_), .A2(new_n594_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n682_), .A2(new_n365_), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n745_), .B2(new_n742_), .ZN(G1336gat));
  INV_X1    g545(.A(G92gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n741_), .A2(new_n747_), .A3(new_n629_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n694_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n682_), .A2(new_n749_), .A3(new_n744_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n750_), .B2(new_n747_), .ZN(G1337gat));
  NOR2_X1   g550(.A1(new_n682_), .A2(new_n744_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n263_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n262_), .A2(new_n459_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n753_), .A2(G99gat), .B1(new_n741_), .B2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g555(.A(new_n460_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n741_), .A2(new_n342_), .A3(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n682_), .A2(new_n343_), .A3(new_n744_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G106gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT111), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n676_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n670_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT107), .B1(new_n764_), .B2(KEYINPUT43), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n679_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n672_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n744_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n342_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n760_), .A4(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n760_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n762_), .B(new_n771_), .C1(new_n772_), .C2(KEYINPUT112), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n774_), .B(new_n760_), .C1(new_n769_), .C2(G106gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n758_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n758_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  INV_X1    g579(.A(G113gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n596_), .B1(new_n576_), .B2(new_n513_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n608_), .B1(new_n599_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n604_), .B2(new_n597_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n553_), .A2(new_n554_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n555_), .B1(new_n787_), .B2(KEYINPUT55), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n553_), .A2(KEYINPUT55), .A3(new_n554_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n564_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT56), .B(new_n564_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n786_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT114), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(KEYINPUT114), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n786_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n622_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n785_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n563_), .A2(new_n610_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n795_), .B2(KEYINPUT113), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n792_), .A2(new_n806_), .A3(new_n794_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n803_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n802_), .B1(new_n808_), .B2(new_n533_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n801_), .A2(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n808_), .A2(new_n802_), .A3(new_n533_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n594_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n569_), .A2(new_n623_), .A3(new_n611_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT54), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n365_), .A2(new_n262_), .A3(new_n629_), .A4(new_n342_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT115), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n819_), .A3(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n610_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n822_), .A2(KEYINPUT59), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(KEYINPUT59), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n817_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n815_), .A2(new_n822_), .A3(KEYINPUT59), .A4(new_n816_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n781_), .B1(new_n610_), .B2(KEYINPUT117), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(KEYINPUT117), .B2(new_n781_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n781_), .A2(new_n821_), .B1(new_n827_), .B2(new_n829_), .ZN(G1340gat));
  AOI21_X1  g629(.A(new_n569_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n818_), .A2(new_n820_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n569_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(KEYINPUT60), .B2(new_n832_), .ZN(new_n835_));
  OAI22_X1  g634(.A1(new_n831_), .A2(new_n832_), .B1(new_n833_), .B2(new_n835_), .ZN(G1341gat));
  AOI21_X1  g635(.A(new_n594_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n837_));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n710_), .A2(new_n838_), .ZN(new_n839_));
  OAI22_X1  g638(.A1(new_n837_), .A2(new_n838_), .B1(new_n833_), .B2(new_n839_), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n818_), .A2(new_n533_), .A3(new_n820_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT118), .B(G134gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n621_), .A2(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n841_), .A2(new_n842_), .B1(new_n827_), .B2(new_n844_), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n263_), .A2(new_n343_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n815_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n749_), .A2(new_n447_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n847_), .A2(new_n611_), .A3(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(new_n286_), .ZN(G1344gat));
  NOR3_X1   g649(.A1(new_n847_), .A2(new_n569_), .A3(new_n848_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n287_), .ZN(G1345gat));
  NOR3_X1   g651(.A1(new_n847_), .A2(new_n594_), .A3(new_n848_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n853_), .B(new_n855_), .ZN(G1346gat));
  NOR2_X1   g655(.A1(new_n847_), .A2(new_n848_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G162gat), .B1(new_n857_), .B2(new_n533_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n763_), .A2(G162gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n857_), .B2(new_n859_), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n749_), .A2(new_n447_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n263_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n342_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n815_), .A2(new_n610_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n203_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n866_), .B2(new_n203_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n242_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(G1348gat));
  AND2_X1   g670(.A1(new_n815_), .A2(new_n865_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n570_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT120), .B(G176gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1349gat));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n710_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n210_), .ZN(new_n877_));
  INV_X1    g676(.A(G183gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n876_), .ZN(G1350gat));
  NAND2_X1  g678(.A1(new_n533_), .A2(new_n213_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT122), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n872_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n815_), .A2(new_n622_), .A3(new_n865_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(new_n884_), .A3(G190gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(G190gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n882_), .B1(new_n885_), .B2(new_n886_), .ZN(G1351gat));
  INV_X1    g686(.A(new_n846_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n861_), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n888_), .B(new_n889_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n610_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT123), .B(G197gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n570_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n594_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT124), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n890_), .A2(new_n896_), .A3(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n815_), .A2(new_n846_), .A3(new_n861_), .A4(new_n898_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n903_));
  INV_X1    g702(.A(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n899_), .A2(new_n901_), .A3(new_n903_), .A4(new_n904_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n890_), .B2(new_n533_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n622_), .A2(G218gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT126), .Z(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n890_), .B2(new_n911_), .ZN(G1355gat));
endmodule


