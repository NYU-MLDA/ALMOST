//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT78), .B(G183gat), .Z(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT22), .B(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(new_n212_), .B2(KEYINPUT25), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT79), .B1(new_n226_), .B2(KEYINPUT26), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(KEYINPUT79), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n223_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231_));
  INV_X1    g030(.A(G169gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n215_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n220_), .B1(new_n230_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G204gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G197gat), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G204gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT89), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n240_), .B2(G204gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n238_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(new_n241_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT21), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n244_), .B1(new_n242_), .B2(KEYINPUT21), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n246_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n237_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n209_), .A2(new_n210_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n216_), .B(new_n219_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n228_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n222_), .A2(new_n217_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(new_n211_), .A3(new_n233_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n254_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n206_), .B1(new_n255_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n254_), .B2(new_n263_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n267_), .B(new_n205_), .C1(new_n254_), .C2(new_n237_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT18), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n202_), .B1(new_n269_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n267_), .B1(new_n237_), .B2(new_n254_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n206_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n273_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT94), .B1(new_n254_), .B2(new_n263_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n253_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n279_), .A2(new_n251_), .B1(new_n245_), .B2(new_n243_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n258_), .A4(new_n262_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n205_), .A2(KEYINPUT20), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n237_), .B2(new_n254_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT95), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n276_), .B(new_n277_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n274_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT96), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n283_), .A2(new_n285_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT95), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(KEYINPUT96), .A3(new_n276_), .A4(new_n277_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n276_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n273_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n290_), .B1(new_n300_), .B2(new_n202_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT102), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI211_X1 g102(.A(KEYINPUT102), .B(new_n290_), .C1(new_n300_), .C2(new_n202_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  INV_X1    g109(.A(G155gat), .ZN(new_n311_));
  INV_X1    g110(.A(G162gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT1), .B1(new_n311_), .B2(new_n312_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n309_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n308_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n313_), .A2(new_n310_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(KEYINPUT84), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT84), .B1(new_n327_), .B2(new_n328_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n318_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT28), .B1(new_n332_), .B2(KEYINPUT29), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n328_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n317_), .B1(new_n336_), .B2(new_n329_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n333_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n333_), .B2(new_n340_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G22gat), .B(G50gat), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n343_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n333_), .A2(new_n340_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT85), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n349_), .B2(new_n342_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT86), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT90), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT88), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n254_), .B2(KEYINPUT87), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n332_), .A2(KEYINPUT29), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n254_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n358_), .B1(new_n359_), .B2(new_n254_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n353_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n254_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n357_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n353_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(KEYINPUT91), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n346_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n349_), .A2(new_n345_), .A3(new_n342_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT91), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n373_), .B(new_n353_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n351_), .A2(new_n368_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n363_), .A3(new_n367_), .A4(new_n371_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(KEYINPUT92), .A3(new_n376_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(G71gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G99gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G15gat), .B(G43gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT82), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n390_), .B(new_n392_), .Z(new_n393_));
  NOR2_X1   g192(.A1(new_n385_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n393_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n383_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G127gat), .B(G134gat), .Z(new_n397_));
  XOR2_X1   g196(.A(G113gat), .B(G120gat), .Z(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OR3_X1    g200(.A1(new_n394_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n399_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n332_), .B2(KEYINPUT97), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT97), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n337_), .A2(new_n407_), .A3(new_n399_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(KEYINPUT98), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(KEYINPUT99), .B(KEYINPUT4), .Z(new_n415_));
  NOR3_X1   g214(.A1(new_n405_), .A2(new_n337_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n409_), .B2(KEYINPUT4), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n414_), .B1(new_n417_), .B2(new_n413_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G1gat), .B(G29gat), .Z(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT100), .B(G85gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G57gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n414_), .B(new_n423_), .C1(new_n417_), .C2(new_n413_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n404_), .A2(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n305_), .A2(new_n381_), .A3(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n375_), .A2(KEYINPUT92), .A3(new_n376_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT92), .B1(new_n375_), .B2(new_n376_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n428_), .B(new_n301_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n277_), .A2(KEYINPUT32), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n294_), .A2(new_n295_), .B1(new_n206_), .B2(new_n275_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(KEYINPUT101), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n265_), .A2(new_n268_), .A3(new_n434_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT101), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n427_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n425_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n418_), .A2(KEYINPUT33), .A3(new_n424_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n417_), .A2(new_n413_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(new_n423_), .C1(new_n413_), .C2(new_n410_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n440_), .B1(new_n446_), .B2(new_n300_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n404_), .B1(new_n433_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n430_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G15gat), .B(G22gat), .ZN(new_n451_));
  INV_X1    g250(.A(G1gat), .ZN(new_n452_));
  INV_X1    g251(.A(G8gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT14), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G8gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n459_), .A2(KEYINPUT69), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(KEYINPUT69), .ZN(new_n461_));
  XOR2_X1   g260(.A(G43gat), .B(G50gat), .Z(new_n462_));
  OR3_X1    g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n462_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT73), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT73), .B1(new_n463_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n458_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT15), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT15), .B1(new_n463_), .B2(new_n464_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n457_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G229gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT74), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT75), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n467_), .A2(new_n470_), .A3(new_n475_), .A4(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n463_), .A2(new_n464_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT73), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT73), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n457_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n467_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n471_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G113gat), .B(G141gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT76), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G169gat), .B(G197gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n474_), .A2(new_n476_), .A3(new_n484_), .A4(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT77), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n473_), .A2(KEYINPUT75), .B1(new_n482_), .B2(new_n483_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(KEYINPUT77), .A3(new_n476_), .A4(new_n488_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n476_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n488_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n450_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n468_), .A2(new_n469_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G85gat), .B(G92gat), .Z(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  INV_X1    g303(.A(G106gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n389_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT7), .ZN(new_n507_));
  AND3_X1   g306(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n504_), .A2(new_n511_), .A3(new_n389_), .A4(new_n505_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n507_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n503_), .B1(new_n513_), .B2(KEYINPUT66), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT10), .B(G99gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n505_), .A2(new_n517_), .B1(new_n503_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n520_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n510_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G85gat), .B(G92gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT66), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n515_), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n519_), .A2(new_n522_), .B1(new_n513_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n516_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT34), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n502_), .A2(new_n527_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(new_n528_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n527_), .A2(new_n477_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G190gat), .B(G218gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G134gat), .B(G162gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT36), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n531_), .A2(new_n528_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n516_), .A2(new_n526_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n535_), .B(new_n542_), .C1(new_n501_), .C2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n533_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT70), .B1(new_n531_), .B2(new_n528_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n539_), .A2(KEYINPUT36), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n536_), .A2(new_n541_), .A3(new_n547_), .A4(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n536_), .A2(new_n547_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n551_), .B2(new_n540_), .ZN(new_n552_));
  AOI211_X1 g351(.A(KEYINPUT71), .B(new_n541_), .C1(new_n536_), .C2(new_n547_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(KEYINPUT37), .B(new_n549_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n457_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(KEYINPUT11), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT67), .ZN(new_n563_));
  INV_X1    g362(.A(G57gat), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(G64gat), .ZN(new_n565_));
  INV_X1    g364(.A(G64gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(G57gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n563_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(G57gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(G64gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(KEYINPUT67), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n562_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n568_), .A2(new_n562_), .A3(new_n571_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n575_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n573_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n569_), .A2(new_n570_), .A3(KEYINPUT67), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT67), .B1(new_n569_), .B2(new_n570_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n581_), .A2(new_n582_), .A3(KEYINPUT11), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT68), .B1(new_n583_), .B2(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n572_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n561_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n595_), .B1(new_n588_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n559_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n578_), .A2(new_n579_), .A3(new_n573_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n572_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n543_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n580_), .A2(new_n586_), .A3(new_n527_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(KEYINPUT12), .A3(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n580_), .A2(new_n586_), .A3(new_n527_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT12), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n603_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n527_), .B1(new_n580_), .B2(new_n586_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n602_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT13), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n612_), .A2(new_n615_), .A3(new_n620_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n623_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n601_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n500_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n452_), .A3(new_n427_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT38), .ZN(new_n632_));
  INV_X1    g431(.A(new_n554_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT103), .B1(new_n450_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n635_), .B(new_n554_), .C1(new_n430_), .C2(new_n449_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n627_), .A2(new_n499_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n599_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(new_n427_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n632_), .B1(new_n642_), .B2(new_n452_), .ZN(G1324gat));
  NAND3_X1  g442(.A1(new_n630_), .A2(new_n453_), .A3(new_n305_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n303_), .A2(new_n304_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n381_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n429_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n433_), .A2(new_n448_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n404_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n635_), .B1(new_n653_), .B2(new_n554_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n636_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n305_), .B(new_n640_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT104), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n637_), .A2(new_n658_), .A3(new_n305_), .A4(new_n640_), .ZN(new_n659_));
  AND4_X1   g458(.A1(new_n645_), .A2(new_n657_), .A3(G8gat), .A4(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n453_), .B1(new_n656_), .B2(KEYINPUT104), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n645_), .B1(new_n661_), .B2(new_n659_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n644_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT40), .B(new_n644_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  NAND3_X1  g466(.A1(new_n637_), .A2(new_n404_), .A3(new_n640_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(KEYINPUT105), .A3(G15gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT105), .B1(new_n668_), .B2(G15gat), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n669_), .A2(new_n670_), .A3(KEYINPUT41), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT41), .B1(new_n669_), .B2(new_n670_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n629_), .A2(G15gat), .A3(new_n651_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT106), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n674_), .ZN(G1326gat));
  INV_X1    g474(.A(new_n641_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G22gat), .B1(new_n676_), .B2(new_n647_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT42), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT42), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n647_), .A2(G22gat), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT107), .Z(new_n681_));
  OAI22_X1  g480(.A1(new_n678_), .A2(new_n679_), .B1(new_n629_), .B2(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n653_), .A2(new_n683_), .A3(new_n558_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n653_), .B2(new_n558_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n639_), .A2(new_n600_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT44), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n688_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(G29gat), .A3(new_n427_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n633_), .A2(new_n599_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n627_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n500_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n428_), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n689_), .A2(new_n691_), .B1(G29gat), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT108), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n694_), .A2(G36gat), .A3(new_n646_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT45), .Z(new_n699_));
  NAND2_X1  g498(.A1(new_n690_), .A2(new_n305_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G36gat), .B1(new_n689_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND3_X1  g505(.A1(new_n690_), .A2(G43gat), .A3(new_n404_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n694_), .A2(new_n651_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n689_), .A2(new_n707_), .B1(G43gat), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g509(.A(new_n694_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G50gat), .B1(new_n711_), .B2(new_n381_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n689_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n690_), .A2(G50gat), .A3(new_n381_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1331gat));
  NOR2_X1   g514(.A1(new_n450_), .A2(new_n498_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n627_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n601_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n564_), .A3(new_n427_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n494_), .A2(new_n497_), .A3(new_n600_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n717_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n637_), .A2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n427_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n722_), .B1(new_n727_), .B2(new_n564_), .ZN(G1332gat));
  NAND3_X1  g527(.A1(new_n721_), .A2(new_n566_), .A3(new_n305_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n726_), .A2(new_n305_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G64gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT48), .B(new_n566_), .C1(new_n726_), .C2(new_n305_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1333gat));
  NAND3_X1  g533(.A1(new_n721_), .A2(new_n387_), .A3(new_n404_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n726_), .A2(new_n404_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G71gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT49), .B(new_n387_), .C1(new_n726_), .C2(new_n404_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n721_), .A2(new_n741_), .A3(new_n381_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n637_), .A2(new_n381_), .A3(new_n725_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(G78gat), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n743_), .A3(G78gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n717_), .A2(new_n692_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n716_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n427_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n717_), .A2(new_n498_), .A3(new_n600_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n754_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT111), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n754_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n427_), .A2(G85gat), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT112), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n753_), .B1(new_n759_), .B2(new_n761_), .ZN(G1336gat));
  NOR3_X1   g561(.A1(new_n751_), .A2(G92gat), .A3(new_n646_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n646_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n765_));
  INV_X1    g564(.A(G92gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n752_), .A2(new_n404_), .A3(new_n517_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n651_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n389_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n752_), .A2(new_n505_), .A3(new_n381_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n381_), .B(new_n754_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G106gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G106gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT114), .B1(new_n627_), .B2(new_n724_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n723_), .A2(new_n625_), .A3(new_n783_), .A4(new_n626_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n781_), .B1(new_n785_), .B2(new_n559_), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT54), .B(new_n558_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n607_), .A2(KEYINPUT12), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n614_), .B2(KEYINPUT12), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT115), .B(new_n789_), .C1(new_n791_), .C2(new_n603_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n612_), .B2(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n612_), .A2(KEYINPUT55), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n603_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n792_), .A2(new_n794_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n620_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n624_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n488_), .B1(new_n482_), .B2(new_n472_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n467_), .A2(new_n470_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n472_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n494_), .A2(new_n804_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n620_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(KEYINPUT116), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT58), .B1(new_n803_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n803_), .A2(KEYINPUT58), .A3(new_n810_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n558_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n498_), .A2(new_n804_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n494_), .B(new_n807_), .C1(new_n622_), .C2(new_n624_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n554_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT57), .B(new_n554_), .C1(new_n816_), .C2(new_n818_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n814_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n788_), .B1(new_n823_), .B2(new_n599_), .ZN(new_n824_));
  NOR4_X1   g623(.A1(new_n305_), .A2(new_n381_), .A3(new_n651_), .A4(new_n428_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n498_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n829_));
  NOR2_X1   g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n786_), .A2(new_n787_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n821_), .A2(new_n822_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n803_), .A2(KEYINPUT58), .A3(new_n810_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n833_), .A2(new_n811_), .A3(new_n559_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n599_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n831_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT118), .B1(new_n823_), .B2(new_n599_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT59), .B1(new_n824_), .B2(new_n826_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n499_), .A2(KEYINPUT119), .ZN(new_n842_));
  MUX2_X1   g641(.A(KEYINPUT119), .B(new_n842_), .S(G113gat), .Z(new_n843_));
  AOI21_X1  g642(.A(new_n828_), .B1(new_n841_), .B2(new_n843_), .ZN(G1340gat));
  NAND3_X1  g643(.A1(new_n839_), .A2(new_n627_), .A3(new_n840_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n839_), .A2(KEYINPUT120), .A3(new_n627_), .A4(new_n840_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(G120gat), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(G120gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n717_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n827_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n850_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(G1341gat));
  NAND4_X1  g652(.A1(new_n839_), .A2(G127gat), .A3(new_n600_), .A4(new_n840_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n835_), .A2(new_n831_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n600_), .A3(new_n825_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n858_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT121), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n854_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT122), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n854_), .A2(new_n861_), .A3(new_n864_), .A4(new_n859_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1342gat));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n827_), .A2(new_n867_), .A3(new_n633_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n841_), .A2(new_n558_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1343gat));
  NOR3_X1   g669(.A1(new_n647_), .A2(new_n428_), .A3(new_n404_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n855_), .A2(new_n646_), .A3(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n499_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n320_), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n717_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n321_), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n872_), .A2(new_n599_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n872_), .B2(new_n559_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n633_), .A2(new_n312_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n872_), .B2(new_n881_), .ZN(G1347gat));
  NAND2_X1  g681(.A1(new_n835_), .A2(new_n836_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n823_), .A2(KEYINPUT118), .A3(new_n599_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n831_), .A3(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n646_), .A2(new_n429_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(new_n381_), .A3(new_n499_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(new_n214_), .A3(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n232_), .B1(new_n885_), .B2(new_n888_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(KEYINPUT62), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n892_), .B(new_n232_), .C1(new_n885_), .C2(new_n888_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT123), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n888_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G169gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n892_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n890_), .A2(KEYINPUT62), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .A4(new_n889_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n894_), .A2(new_n900_), .ZN(G1348gat));
  NAND2_X1  g700(.A1(new_n855_), .A2(new_n647_), .ZN(new_n902_));
  NOR4_X1   g701(.A1(new_n902_), .A2(new_n215_), .A3(new_n717_), .A4(new_n887_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n887_), .A2(new_n381_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n885_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n627_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n906_), .B2(new_n215_), .ZN(G1349gat));
  NOR2_X1   g706(.A1(new_n599_), .A2(new_n259_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n885_), .A2(new_n904_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n902_), .A2(new_n599_), .A3(new_n887_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n212_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n909_), .A2(new_n910_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(G1350gat));
  NAND3_X1  g714(.A1(new_n905_), .A2(new_n228_), .A3(new_n633_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n905_), .A2(new_n558_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n918_), .B2(new_n226_), .ZN(G1351gat));
  NAND3_X1  g718(.A1(new_n381_), .A2(new_n651_), .A3(new_n428_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT125), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n305_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n824_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n498_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n627_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g726(.A(new_n923_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT63), .B(G211gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n928_), .A2(new_n599_), .A3(new_n929_), .ZN(new_n930_));
  AOI211_X1 g729(.A(KEYINPUT63), .B(G211gat), .C1(new_n923_), .C2(new_n600_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1354gat));
  NAND2_X1  g731(.A1(new_n558_), .A2(G218gat), .ZN(new_n933_));
  XOR2_X1   g732(.A(new_n933_), .B(KEYINPUT126), .Z(new_n934_));
  NOR2_X1   g733(.A1(new_n928_), .A2(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G218gat), .B1(new_n923_), .B2(new_n633_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937_));
  OR3_X1    g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1355gat));
endmodule


