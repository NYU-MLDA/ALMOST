//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  AOI21_X1  g000(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND3_X1  g002(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT66), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n206_));
  INV_X1    g005(.A(new_n204_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT10), .B(G99gat), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n209_), .A2(new_n211_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n207_), .A2(new_n202_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n213_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT67), .A3(new_n220_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n218_), .B1(new_n229_), .B2(new_n215_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n215_), .A2(new_n218_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n221_), .A2(new_n222_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n209_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n217_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G78gat), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n234_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT12), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n241_), .B(new_n217_), .C1(new_n230_), .C2(new_n233_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(KEYINPUT12), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT64), .Z(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT65), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n245_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(G204gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT5), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n255_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n252_), .A2(new_n254_), .A3(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(KEYINPUT13), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(KEYINPUT13), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT69), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT15), .ZN(new_n272_));
  INV_X1    g071(.A(G29gat), .ZN(new_n273_));
  INV_X1    g072(.A(G36gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G43gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G29gat), .A2(G36gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G50gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n276_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G29gat), .B(G36gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G43gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(G50gat), .B1(new_n284_), .B2(new_n278_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n272_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n280_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(G50gat), .A3(new_n278_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT15), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n234_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n282_), .A2(new_n285_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(new_n217_), .C1(new_n230_), .C2(new_n233_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT34), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n234_), .A2(new_n290_), .A3(KEYINPUT71), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n293_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n298_), .A2(new_n300_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n304_), .A2(KEYINPUT72), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT72), .B1(new_n304_), .B2(new_n305_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n305_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n293_), .A2(new_n302_), .A3(new_n309_), .A4(new_n303_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT74), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n271_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G190gat), .B(G218gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G134gat), .ZN(new_n314_));
  INV_X1    g113(.A(G162gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT36), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n304_), .A2(new_n305_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n304_), .A2(KEYINPUT72), .A3(new_n305_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n310_), .B(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT75), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n312_), .A2(new_n317_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n324_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT36), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n316_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT73), .Z(new_n330_));
  OR2_X1    g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT37), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n327_), .A2(new_n330_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n317_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n335_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G15gat), .B(G22gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G1gat), .A2(G8gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT14), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G8gat), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n345_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G231gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(new_n242_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT16), .B(G183gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G211gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G155gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT17), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n351_), .B2(KEYINPUT76), .ZN(new_n358_));
  MUX2_X1   g157(.A(new_n357_), .B(KEYINPUT17), .S(new_n358_), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n340_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n270_), .A2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n362_), .A2(KEYINPUT77), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT2), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT91), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT89), .B(KEYINPUT3), .ZN(new_n371_));
  NOR2_X1   g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n374_));
  NOR2_X1   g173(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n370_), .B(new_n372_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n367_), .B(new_n369_), .C1(new_n373_), .C2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G155gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n315_), .A3(KEYINPUT87), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(G155gat), .B2(G162gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT92), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n380_), .A2(new_n382_), .A3(new_n386_), .A4(new_n383_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT88), .B1(new_n383_), .B2(KEYINPUT1), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(G155gat), .A4(G162gat), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n383_), .A2(KEYINPUT1), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n380_), .A2(new_n396_), .A3(new_n382_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n372_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n366_), .ZN(new_n399_));
  AND4_X1   g198(.A1(KEYINPUT93), .A2(new_n389_), .A3(new_n390_), .A4(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n378_), .A2(new_n388_), .B1(new_n398_), .B2(new_n366_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT93), .B1(new_n401_), .B2(new_n390_), .ZN(new_n402_));
  OAI21_X1  g201(.A(G22gat), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n389_), .A2(new_n390_), .A3(new_n399_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G22gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(KEYINPUT93), .A3(new_n390_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n403_), .A2(G50gat), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(G50gat), .B1(new_n403_), .B2(new_n409_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n365_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n390_), .B1(new_n389_), .B2(new_n399_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G211gat), .B(G218gat), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n257_), .A2(G197gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n257_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n420_));
  INV_X1    g219(.A(G197gat), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n419_), .A2(new_n420_), .B1(new_n421_), .B2(G204gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT21), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n416_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  OR3_X1    g223(.A1(new_n257_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT95), .B1(new_n257_), .B2(G197gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n417_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT21), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n422_), .A2(new_n423_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n416_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n414_), .B1(new_n415_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n431_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n434_), .B(new_n413_), .C1(new_n401_), .C2(new_n390_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n436_), .A2(KEYINPUT98), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n400_), .A2(new_n402_), .A3(G22gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n407_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n280_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n403_), .A2(G50gat), .A3(new_n409_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n364_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n412_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n433_), .A2(KEYINPUT98), .A3(new_n435_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT97), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT97), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n433_), .A2(new_n446_), .A3(KEYINPUT98), .A4(new_n435_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G78gat), .B(G106gat), .Z(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n451_), .A3(new_n447_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n443_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n443_), .A2(new_n453_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT23), .ZN(new_n459_));
  OR2_X1    g258(.A1(G183gat), .A2(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT22), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n260_), .B1(new_n462_), .B2(KEYINPUT85), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G169gat), .ZN(new_n464_));
  INV_X1    g263(.A(G169gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n260_), .C1(new_n462_), .C2(KEYINPUT85), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G183gat), .A2(G190gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT84), .B1(new_n468_), .B2(KEYINPUT83), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT23), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n469_), .A2(new_n470_), .B1(KEYINPUT84), .B2(new_n468_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT25), .B(G183gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT26), .B(G190gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n465_), .A2(new_n260_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G169gat), .A2(G176gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT24), .A3(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n476_), .B(new_n479_), .C1(KEYINPUT24), .C2(new_n477_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n467_), .B1(new_n473_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT30), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n467_), .B(new_n483_), .C1(new_n473_), .C2(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT86), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G127gat), .B(G134gat), .ZN(new_n487_));
  INV_X1    g286(.A(G113gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G120gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n482_), .A2(new_n492_), .A3(new_n484_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G71gat), .B(G99gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(G15gat), .B(G43gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G227gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n491_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(new_n491_), .A3(new_n498_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n490_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  INV_X1    g302(.A(G120gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n489_), .B(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n503_), .A2(new_n505_), .A3(new_n499_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n486_), .B1(new_n502_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n503_), .B2(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(new_n490_), .A3(new_n501_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT86), .A4(new_n485_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G64gat), .B(G92gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(G36gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT100), .B(G8gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n434_), .A2(new_n481_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n459_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n480_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n460_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n478_), .B1(new_n473_), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G169gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(G176gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n521_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n519_), .B(KEYINPUT20), .C1(new_n527_), .C2(new_n434_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G226gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT19), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT20), .ZN(new_n533_));
  INV_X1    g332(.A(new_n481_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n432_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n434_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n530_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT104), .B1(new_n532_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n528_), .A2(new_n530_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n531_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(KEYINPUT32), .B(new_n518_), .C1(new_n538_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n518_), .A2(KEYINPUT32), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n532_), .A2(new_n537_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(KEYINPUT104), .ZN(new_n545_));
  XOR2_X1   g344(.A(G1gat), .B(G29gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G57gat), .B(G85gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n401_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n490_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n505_), .A2(new_n401_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT4), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n505_), .A2(new_n401_), .A3(KEYINPUT4), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G225gat), .A2(G233gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT101), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n550_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n550_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n542_), .B(new_n545_), .C1(new_n561_), .C2(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n532_), .A2(new_n537_), .A3(new_n517_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n517_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT103), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n559_), .A2(new_n560_), .A3(new_n550_), .A4(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n554_), .A2(new_n556_), .A3(new_n555_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n552_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n563_), .A3(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n568_), .A2(new_n570_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n565_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n457_), .A2(new_n511_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n567_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT105), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT27), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n541_), .B2(new_n517_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(KEYINPUT105), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n581_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n564_), .A2(new_n561_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n582_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n507_), .A2(new_n510_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n454_), .A2(new_n455_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n452_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n451_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n594_), .A2(new_n437_), .A3(new_n442_), .A4(new_n412_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n443_), .A2(new_n453_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n511_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n589_), .B1(new_n591_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n579_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT79), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n287_), .A2(new_n288_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n348_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n346_), .A2(new_n287_), .A3(new_n347_), .A4(new_n288_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(KEYINPUT78), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n348_), .A2(new_n601_), .A3(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n604_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n286_), .A2(new_n289_), .B1(new_n347_), .B2(new_n346_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n603_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n610_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n600_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G113gat), .B(G141gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(G197gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT80), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(G169gat), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT80), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n615_), .B(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n465_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT81), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n617_), .A2(new_n620_), .A3(KEYINPUT81), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n610_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n605_), .A3(new_n603_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n604_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(KEYINPUT79), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n613_), .A2(new_n625_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT82), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n628_), .A3(new_n621_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT82), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n613_), .A2(new_n625_), .A3(new_n629_), .A4(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n362_), .B2(KEYINPUT77), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n363_), .A2(new_n599_), .A3(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G1gat), .A3(new_n586_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n360_), .B1(new_n579_), .B2(new_n598_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(new_n332_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n269_), .A2(new_n636_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n586_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n645_), .A3(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n585_), .A2(new_n587_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n642_), .A2(new_n643_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(G8gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n650_), .B2(G8gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n648_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(G8gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT106), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(KEYINPUT39), .A3(new_n652_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n363_), .A2(new_n599_), .A3(new_n637_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n649_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(G8gat), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n655_), .A2(new_n658_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n655_), .A2(new_n662_), .A3(new_n658_), .A4(KEYINPUT40), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  INV_X1    g466(.A(new_n644_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n590_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G15gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT107), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n672_), .A3(G15gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n638_), .A2(G15gat), .A3(new_n511_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(KEYINPUT41), .A3(new_n673_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(G1326gat));
  AND2_X1   g478(.A1(new_n456_), .A2(KEYINPUT108), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n456_), .A2(KEYINPUT108), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n659_), .A2(new_n407_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n682_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G22gat), .B1(new_n644_), .B2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n340_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n590_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n595_), .A2(new_n511_), .A3(new_n596_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n588_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  AOI221_X4 g493(.A(new_n590_), .B1(new_n565_), .B2(new_n577_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n340_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  OAI221_X1 g496(.A(new_n340_), .B1(new_n690_), .B2(new_n689_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n643_), .A4(new_n360_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n586_), .A2(new_n273_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n643_), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n702_), .B(new_n359_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n703_), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n699_), .A2(new_n643_), .A3(new_n360_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n700_), .B(new_n701_), .C1(new_n704_), .C2(new_n708_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n332_), .B(new_n359_), .C1(new_n579_), .C2(new_n598_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n643_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n273_), .B1(new_n711_), .B2(new_n586_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(KEYINPUT111), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1328gat));
  NAND4_X1  g516(.A1(new_n710_), .A2(new_n274_), .A3(new_n643_), .A4(new_n649_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT45), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n700_), .A2(new_n649_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT110), .B1(new_n703_), .B2(KEYINPUT44), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n706_), .A2(new_n705_), .A3(new_n707_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n723_), .B2(new_n274_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT46), .B(new_n719_), .C1(new_n723_), .C2(new_n274_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NOR2_X1   g527(.A1(new_n511_), .A2(new_n276_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n700_), .B(new_n729_), .C1(new_n704_), .C2(new_n708_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n276_), .B1(new_n711_), .B2(new_n511_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT47), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(new_n734_), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1330gat));
  AOI22_X1  g535(.A1(new_n721_), .A2(new_n722_), .B1(KEYINPUT44), .B2(new_n703_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n457_), .A2(new_n280_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n710_), .A2(new_n643_), .A3(new_n682_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n737_), .A2(new_n738_), .B1(new_n280_), .B2(new_n739_), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n270_), .A2(new_n635_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n642_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n586_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n340_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n269_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n635_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n641_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n586_), .B1(new_n749_), .B2(KEYINPUT112), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(KEYINPUT112), .B2(new_n749_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n744_), .B1(new_n751_), .B2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n742_), .B2(new_n660_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(KEYINPUT113), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(KEYINPUT113), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(KEYINPUT48), .A3(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n749_), .A2(new_n649_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n758_), .B(new_n759_), .C1(G64gat), .C2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n742_), .B2(new_n511_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT49), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT49), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n511_), .A2(G71gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT114), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n763_), .A2(new_n764_), .B1(new_n748_), .B2(new_n766_), .ZN(G1334gat));
  OR3_X1    g566(.A1(new_n748_), .A2(G78gat), .A3(new_n684_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G78gat), .B1(new_n742_), .B2(new_n684_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  AND2_X1   g571(.A1(new_n741_), .A2(new_n710_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n586_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G85gat), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n360_), .B(new_n747_), .C1(new_n699_), .C2(KEYINPUT115), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n776_), .A2(new_n586_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n775_), .B1(new_n779_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g579(.A(G92gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n773_), .A2(new_n781_), .A3(new_n649_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n776_), .A2(new_n778_), .A3(new_n660_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n781_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT116), .ZN(G1337gat));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT51), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT118), .Z(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n773_), .A2(new_n212_), .A3(new_n590_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n747_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n699_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n777_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n778_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n590_), .A3(new_n360_), .A4(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n790_), .B1(new_n795_), .B2(G99gat), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n786_), .A2(KEYINPUT51), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n789_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n797_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n776_), .A2(new_n778_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n226_), .B1(new_n800_), .B2(new_n590_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n799_), .B(new_n788_), .C1(new_n801_), .C2(new_n790_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(new_n802_), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n773_), .A2(new_n456_), .A3(new_n213_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n699_), .A2(new_n456_), .A3(new_n360_), .A4(new_n747_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(G106gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(G106gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n247_), .A2(new_n251_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n252_), .A2(KEYINPUT55), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n247_), .A2(new_n814_), .A3(new_n251_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n812_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n262_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n811_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n819_));
  AOI211_X1 g618(.A(KEYINPUT55), .B(new_n250_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n819_), .A2(new_n820_), .B1(new_n251_), .B2(new_n247_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n262_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n626_), .A2(new_n606_), .A3(new_n603_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n604_), .A2(new_n605_), .A3(new_n608_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n824_), .A2(new_n617_), .A3(new_n825_), .A4(new_n620_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n826_), .A2(new_n632_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(new_n264_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n264_), .A4(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n340_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n635_), .A2(new_n264_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n822_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n262_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n265_), .A2(new_n827_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n332_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n838_), .B2(new_n332_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n832_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT119), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n832_), .B(new_n844_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n360_), .A3(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n361_), .A2(new_n746_), .A3(new_n636_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT54), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n361_), .A2(new_n849_), .A3(new_n746_), .A4(new_n636_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n846_), .A2(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n692_), .A2(new_n586_), .A3(new_n649_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n488_), .B1(new_n854_), .B2(new_n636_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n842_), .A2(new_n360_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT121), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n842_), .A2(new_n861_), .A3(new_n360_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n851_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n853_), .A3(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n858_), .A2(G113gat), .A3(new_n635_), .A4(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT120), .B(new_n488_), .C1(new_n854_), .C2(new_n636_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n857_), .A2(new_n866_), .A3(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(new_n854_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n504_), .B1(new_n746_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n869_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n504_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n865_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n864_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n270_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n871_), .B1(new_n874_), .B2(new_n504_), .ZN(G1341gat));
  AOI21_X1  g674(.A(G127gat), .B1(new_n869_), .B2(new_n359_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n858_), .A2(G127gat), .A3(new_n865_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n359_), .ZN(G1342gat));
  INV_X1    g677(.A(new_n332_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G134gat), .B1(new_n869_), .B2(new_n879_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n872_), .A2(new_n873_), .A3(new_n745_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g681(.A(new_n693_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n649_), .A2(new_n586_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n635_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g685(.A(new_n270_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n883_), .A2(new_n887_), .A3(new_n884_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n883_), .A2(new_n884_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n360_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT61), .B(G155gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  NOR3_X1   g692(.A1(new_n890_), .A2(new_n315_), .A3(new_n745_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n883_), .A2(new_n879_), .A3(new_n884_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n315_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(KEYINPUT122), .A3(new_n315_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n894_), .B1(new_n898_), .B2(new_n899_), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n660_), .A2(new_n774_), .A3(new_n511_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n684_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n863_), .A2(new_n635_), .A3(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n903_), .A2(G169gat), .A3(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n904_), .A2(new_n905_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n908_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n903_), .A2(G169gat), .A3(new_n910_), .A4(new_n906_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n909_), .B(new_n911_), .C1(new_n525_), .C2(new_n903_), .ZN(G1348gat));
  NAND2_X1  g711(.A1(new_n863_), .A2(new_n902_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n260_), .B1(new_n913_), .B2(new_n746_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n456_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n915_), .A2(G176gat), .A3(new_n887_), .A4(new_n901_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1349gat));
  NAND4_X1  g716(.A1(new_n852_), .A2(new_n457_), .A3(new_n359_), .A4(new_n901_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(G183gat), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n915_), .A2(KEYINPUT125), .A3(new_n359_), .A4(new_n901_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n913_), .A2(new_n474_), .A3(new_n360_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n913_), .B2(new_n745_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n879_), .A2(new_n475_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n913_), .B2(new_n927_), .ZN(G1351gat));
  NOR2_X1   g727(.A1(new_n693_), .A2(new_n774_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(KEYINPUT126), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n660_), .B1(new_n929_), .B2(KEYINPUT126), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n635_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G197gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n933_), .A2(new_n421_), .A3(new_n635_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1352gat));
  NAND3_X1  g736(.A1(new_n931_), .A2(new_n887_), .A3(new_n932_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n931_), .A2(new_n359_), .A3(new_n932_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT63), .B(G211gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n940_), .B2(new_n943_), .ZN(G1354gat));
  XOR2_X1   g743(.A(KEYINPUT127), .B(G218gat), .Z(new_n945_));
  AOI21_X1  g744(.A(new_n945_), .B1(new_n933_), .B2(new_n879_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n340_), .A2(new_n945_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n933_), .B2(new_n947_), .ZN(G1355gat));
endmodule


