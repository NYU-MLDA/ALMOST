//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT67), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT74), .Z(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT71), .B(G15gat), .Z(new_n207_));
  INV_X1    g006(.A(G22gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209_));
  AND2_X1   g008(.A1(G1gat), .A2(G8gat), .ZN(new_n210_));
  OAI22_X1  g009(.A1(new_n207_), .A2(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(new_n208_), .B2(new_n207_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G1gat), .A2(G8gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n212_), .B(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n206_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n205_), .B(KEYINPUT15), .Z(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n206_), .B(new_n215_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n219_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G169gat), .B(G197gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT75), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n228_), .B(KEYINPUT76), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n224_), .B(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(G127gat), .A2(G134gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G127gat), .A2(G134gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G113gat), .ZN(new_n234_));
  INV_X1    g033(.A(G120gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G113gat), .A2(G120gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT83), .B1(new_n233_), .B2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G127gat), .A2(G134gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n232_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n237_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G113gat), .A2(G120gat), .ZN(new_n243_));
  OAI22_X1  g042(.A1(new_n240_), .A2(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n231_), .A2(new_n236_), .A3(new_n232_), .A4(new_n237_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n239_), .B1(new_n246_), .B2(KEYINPUT83), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT31), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT85), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(G169gat), .B2(G176gat), .ZN(new_n254_));
  INV_X1    g053(.A(G169gat), .ZN(new_n255_));
  INV_X1    g054(.A(G176gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT79), .B(G183gat), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n262_));
  OR3_X1    g061(.A1(new_n262_), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G190gat), .ZN(new_n264_));
  INV_X1    g063(.A(G183gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT25), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT77), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n261_), .A2(new_n263_), .A3(new_n264_), .A4(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT78), .B(KEYINPUT25), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT79), .B1(new_n269_), .B2(G183gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n258_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT80), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n273_), .B(new_n258_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n275_));
  INV_X1    g074(.A(G190gat), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n265_), .A2(new_n276_), .A3(KEYINPUT23), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT23), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n275_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n256_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n279_), .A2(new_n289_), .A3(KEYINPUT23), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n279_), .B2(KEYINPUT23), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n278_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n286_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n282_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT82), .B(G15gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n281_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n271_), .B2(KEYINPUT80), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n294_), .B1(new_n302_), .B2(new_n274_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT30), .B(G43gat), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G71gat), .B(G99gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n307_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n300_), .A2(new_n310_), .A3(new_n305_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n248_), .A2(new_n249_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n309_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n252_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n311_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(new_n313_), .A3(new_n312_), .A4(new_n251_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT94), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G155gat), .B(G162gat), .Z(new_n327_));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328_));
  INV_X1    g127(.A(G141gat), .ZN(new_n329_));
  INV_X1    g128(.A(G148gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT86), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(KEYINPUT2), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n331_), .B(new_n332_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT86), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(KEYINPUT2), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n338_), .A2(new_n339_), .B1(G141gat), .B2(G148gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n327_), .B1(new_n336_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G155gat), .ZN(new_n342_));
  INV_X1    g141(.A(G162gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT1), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(G155gat), .A3(G162gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n344_), .B(new_n346_), .C1(G155gat), .C2(G162gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(G141gat), .B(G148gat), .Z(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n326_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n341_), .A2(new_n349_), .A3(new_n352_), .A4(new_n325_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G22gat), .B(G50gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(new_n357_), .A3(new_n353_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT90), .ZN(new_n360_));
  INV_X1    g159(.A(G204gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(G197gat), .ZN(new_n362_));
  INV_X1    g161(.A(G197gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT88), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(G204gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n361_), .A2(KEYINPUT88), .ZN(new_n368_));
  OAI21_X1  g167(.A(G197gat), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n361_), .A2(KEYINPUT88), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(G204gat), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n363_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n362_), .A2(new_n364_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT91), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n371_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n371_), .A2(new_n376_), .A3(KEYINPUT92), .A4(new_n379_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n374_), .A2(new_n375_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n378_), .ZN(new_n385_));
  AOI21_X1  g184(.A(G197gat), .B1(new_n372_), .B2(new_n373_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n378_), .B1(G197gat), .B2(G204gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT89), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n372_), .A2(new_n373_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n363_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n387_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n385_), .A2(new_n377_), .A3(new_n389_), .A4(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n382_), .A2(new_n383_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G228gat), .ZN(new_n396_));
  INV_X1    g195(.A(G233gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n350_), .A2(KEYINPUT29), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n395_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n395_), .B2(new_n400_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT93), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT93), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n395_), .A2(new_n400_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n398_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n395_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n359_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n359_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n324_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT93), .B1(new_n401_), .B2(new_n402_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n414_), .B2(new_n410_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n401_), .A2(new_n402_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n359_), .B1(new_n416_), .B2(new_n404_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n415_), .A2(new_n417_), .A3(new_n323_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  INV_X1    g219(.A(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT0), .B(G57gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n350_), .A2(new_n247_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n341_), .A2(new_n349_), .A3(new_n246_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT4), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT4), .B1(new_n350_), .B2(new_n247_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n426_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT98), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT98), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n427_), .A2(new_n436_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n425_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n441_));
  OAI211_X1 g240(.A(G225gat), .B(G233gat), .C1(new_n441_), .C2(new_n431_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(new_n424_), .A3(new_n437_), .A4(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G8gat), .B(G36gat), .ZN(new_n446_));
  INV_X1    g245(.A(G92gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT18), .B(G64gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n382_), .A2(new_n383_), .A3(new_n394_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT20), .B1(new_n303_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n275_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n276_), .A2(KEYINPUT26), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT26), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n262_), .A2(G183gat), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n266_), .A2(new_n459_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n280_), .A2(KEYINPUT81), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n277_), .B1(new_n465_), .B2(new_n290_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n457_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n293_), .A2(KEYINPUT96), .A3(new_n463_), .A4(new_n458_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n278_), .A2(new_n280_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n286_), .B1(new_n288_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n456_), .B1(new_n395_), .B2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n453_), .A2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n393_), .A2(new_n389_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n377_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n384_), .B2(new_n378_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n476_), .A2(new_n478_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n282_), .A2(new_n479_), .A3(new_n383_), .A4(new_n295_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(new_n395_), .B2(new_n473_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n456_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n451_), .B1(new_n475_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n482_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n456_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n471_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n486_), .B1(new_n452_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n296_), .A2(new_n395_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT20), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n491_), .A3(new_n450_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT97), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n484_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n487_), .A2(new_n491_), .A3(KEYINPUT97), .A4(new_n450_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n464_), .A2(new_n466_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n471_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n499_), .A2(new_n382_), .A3(new_n383_), .A4(new_n394_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT20), .B(new_n500_), .C1(new_n303_), .C2(new_n452_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT99), .A3(new_n486_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n480_), .A2(new_n482_), .A3(new_n456_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT99), .B1(new_n501_), .B2(new_n486_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n451_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(KEYINPUT27), .A3(new_n492_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n419_), .A2(new_n445_), .A3(new_n497_), .A4(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n409_), .A2(new_n324_), .A3(new_n412_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n323_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT33), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n443_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n438_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n514_), .A2(KEYINPUT33), .A3(new_n424_), .A4(new_n442_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n426_), .B1(new_n441_), .B2(new_n431_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(new_n425_), .C1(new_n426_), .C2(new_n429_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n450_), .A2(KEYINPUT32), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n487_), .A2(new_n491_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n444_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n501_), .A2(new_n486_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n503_), .A3(new_n502_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n522_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n511_), .B1(new_n519_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n321_), .B1(new_n508_), .B2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n507_), .A2(new_n497_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n316_), .A2(new_n320_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n532_), .A2(new_n419_), .A3(new_n444_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n530_), .A2(KEYINPUT101), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n508_), .A2(new_n529_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n532_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT101), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n230_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT102), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G71gat), .B(G78gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(G57gat), .B(G64gat), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n543_), .B2(KEYINPUT11), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(KEYINPUT11), .B2(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n541_), .A3(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n215_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G127gat), .B(G155gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT73), .B1(new_n553_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n553_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n558_), .B(KEYINPUT17), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  MUX2_X1   g363(.A(KEYINPUT73), .B(new_n561_), .S(new_n564_), .Z(new_n565_));
  XOR2_X1   g364(.A(G134gat), .B(G162gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT68), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT36), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G85gat), .B(G92gat), .Z(new_n572_));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT6), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT65), .ZN(new_n577_));
  NOR2_X1   g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT7), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n574_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n576_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n573_), .B1(new_n581_), .B2(new_n572_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n572_), .A2(KEYINPUT9), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n421_), .A2(new_n447_), .A3(KEYINPUT9), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT10), .B(G99gat), .Z(new_n586_));
  INV_X1    g385(.A(G106gat), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n577_), .A2(new_n584_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(new_n205_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT66), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n589_), .B(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n583_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n217_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n591_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n598_), .A2(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n591_), .A2(new_n595_), .A3(new_n604_), .A4(new_n600_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n571_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n569_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT69), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT70), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n603_), .A2(new_n605_), .A3(KEYINPUT70), .A4(new_n609_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n606_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n565_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n590_), .A2(new_n548_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n594_), .A2(KEYINPUT12), .A3(new_n548_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n583_), .A2(new_n547_), .A3(new_n589_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT64), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n623_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n626_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(new_n361_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT5), .B(G176gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n633_), .B(new_n634_), .Z(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n631_), .A2(new_n636_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT13), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT13), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n540_), .A2(new_n618_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n646_), .A2(G1gat), .A3(new_n445_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n644_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n565_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n614_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n539_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n445_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n647_), .A2(new_n648_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n649_), .A2(new_n654_), .A3(new_n655_), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n531_), .A2(G8gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n645_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT103), .ZN(new_n659_));
  OAI21_X1  g458(.A(G8gat), .B1(new_n653_), .B2(new_n531_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT39), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n662_), .B(new_n664_), .ZN(G1325gat));
  OAI21_X1  g464(.A(G15gat), .B1(new_n653_), .B2(new_n532_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT41), .Z(new_n667_));
  OR2_X1    g466(.A1(new_n532_), .A2(G15gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n646_), .B2(new_n668_), .ZN(G1326gat));
  NAND3_X1  g468(.A1(new_n645_), .A2(new_n208_), .A3(new_n419_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G22gat), .B1(new_n653_), .B2(new_n511_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n540_), .A2(new_n644_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n614_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n565_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n444_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n616_), .A2(new_n617_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n535_), .A2(KEYINPUT101), .A3(new_n532_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n533_), .A2(new_n531_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n530_), .A2(KEYINPUT101), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n534_), .A2(new_n538_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(new_n686_), .A3(KEYINPUT43), .A4(new_n680_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n644_), .A2(new_n230_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n690_), .A2(new_n651_), .A3(new_n692_), .A4(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(KEYINPUT106), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT106), .B1(new_n694_), .B2(new_n695_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n694_), .A2(new_n695_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(G29gat), .A3(new_n444_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n679_), .B1(new_n699_), .B2(new_n701_), .ZN(G1328gat));
  NOR2_X1   g501(.A1(new_n531_), .A2(G36gat), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OR3_X1    g503(.A1(new_n677_), .A2(KEYINPUT45), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT45), .B1(new_n677_), .B2(new_n704_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n531_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n694_), .A2(new_n695_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n694_), .A2(KEYINPUT106), .A3(new_n695_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n714_), .A2(KEYINPUT107), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n708_), .B(new_n700_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G36gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n707_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT46), .B(new_n707_), .C1(new_n716_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  NOR2_X1   g523(.A1(new_n677_), .A2(new_n532_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n700_), .A2(G43gat), .A3(new_n321_), .ZN(new_n726_));
  OAI22_X1  g525(.A1(G43gat), .A2(new_n725_), .B1(new_n698_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g527(.A1(new_n677_), .A2(G50gat), .A3(new_n511_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n700_), .A2(new_n419_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G50gat), .B1(new_n698_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n732_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1331gat));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  INV_X1    g535(.A(new_n230_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n650_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n691_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n680_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n565_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n741_), .B2(new_n445_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n652_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n444_), .A2(G57gat), .ZN(new_n744_));
  OAI22_X1  g543(.A1(new_n742_), .A2(KEYINPUT109), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(KEYINPUT109), .B2(new_n742_), .ZN(G1332gat));
  OAI21_X1  g545(.A(G64gat), .B1(new_n743_), .B2(new_n531_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT48), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n531_), .A2(G64gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n741_), .B2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT110), .Z(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n743_), .B2(new_n532_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n532_), .A2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n741_), .B2(new_n755_), .ZN(G1334gat));
  OAI21_X1  g555(.A(G78gat), .B1(new_n743_), .B2(new_n511_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n511_), .A2(G78gat), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT112), .Z(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n741_), .B2(new_n760_), .ZN(G1335gat));
  AND2_X1   g560(.A1(new_n692_), .A2(new_n651_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n690_), .A3(new_n738_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n763_), .A2(new_n421_), .A3(new_n445_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n739_), .A2(new_n676_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n444_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1336gat));
  NOR3_X1   g566(.A1(new_n763_), .A2(new_n447_), .A3(new_n531_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G92gat), .B1(new_n765_), .B2(new_n708_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n763_), .B2(new_n532_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n586_), .A3(new_n321_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT113), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n775_), .A2(new_n778_), .B1(new_n776_), .B2(new_n774_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n780_), .ZN(G1338gat));
  OAI21_X1  g582(.A(G106gat), .B1(new_n763_), .B2(new_n511_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT52), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n765_), .A2(new_n587_), .A3(new_n419_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT115), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n788_), .B(new_n790_), .ZN(G1339gat));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n641_), .A2(new_n643_), .A3(new_n230_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n792_), .B(KEYINPUT54), .C1(new_n793_), .C2(new_n618_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n793_), .A2(new_n618_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(KEYINPUT54), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(KEYINPUT54), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n624_), .A2(KEYINPUT55), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n629_), .B2(KEYINPUT118), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n627_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n624_), .A2(new_n801_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n635_), .B1(new_n805_), .B2(KEYINPUT119), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n803_), .A2(new_n807_), .A3(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n808_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n809_), .A2(KEYINPUT120), .A3(new_n810_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n218_), .A2(new_n219_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n221_), .A2(new_n222_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n227_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n227_), .B2(new_n224_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n639_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n814_), .A2(new_n815_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n815_), .A4(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n680_), .A3(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n230_), .A2(new_n639_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n640_), .A2(new_n819_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n675_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT57), .B(new_n675_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n798_), .B1(new_n833_), .B2(new_n651_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n532_), .A2(new_n419_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n708_), .A2(new_n445_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n834_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n737_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n833_), .A2(new_n651_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n798_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n838_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n844_), .B2(new_n835_), .ZN(new_n845_));
  NOR4_X1   g644(.A1(new_n834_), .A2(KEYINPUT59), .A3(new_n836_), .A4(new_n838_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n230_), .A2(new_n234_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n840_), .B1(new_n847_), .B2(new_n848_), .ZN(G1340gat));
  NOR2_X1   g648(.A1(new_n235_), .A2(KEYINPUT60), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n235_), .B1(new_n650_), .B2(KEYINPUT60), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(KEYINPUT121), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n839_), .B(new_n852_), .C1(KEYINPUT121), .C2(new_n851_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n845_), .A2(new_n846_), .A3(new_n650_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n235_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n839_), .B2(new_n565_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT122), .B(G127gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n565_), .A2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT123), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n847_), .B2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n839_), .B2(new_n614_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n680_), .A2(G134gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n847_), .B2(new_n862_), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n321_), .A2(new_n511_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n844_), .A2(new_n737_), .A3(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g665(.A1(new_n844_), .A2(new_n644_), .A3(new_n864_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g667(.A1(new_n844_), .A2(new_n565_), .A3(new_n864_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  INV_X1    g671(.A(new_n864_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n834_), .A2(new_n675_), .A3(new_n838_), .A4(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n874_), .B2(G162gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n844_), .A2(new_n614_), .A3(new_n864_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(KEYINPUT124), .A3(new_n343_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n844_), .A2(G162gat), .A3(new_n680_), .A4(new_n864_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n875_), .A2(new_n877_), .A3(new_n878_), .ZN(G1347gat));
  INV_X1    g678(.A(new_n533_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n834_), .A2(new_n531_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT62), .B(G169gat), .C1(new_n882_), .C2(new_n230_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n834_), .A2(new_n230_), .A3(new_n531_), .A4(new_n880_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n255_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n283_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n883_), .A2(new_n886_), .A3(new_n887_), .ZN(G1348gat));
  NAND2_X1  g687(.A1(new_n881_), .A2(new_n644_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g689(.A(G183gat), .B1(new_n882_), .B2(new_n651_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n881_), .A2(new_n565_), .A3(new_n266_), .A4(new_n462_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1350gat));
  NAND2_X1  g692(.A1(new_n842_), .A2(new_n843_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n614_), .A2(new_n264_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT125), .Z(new_n896_));
  NAND4_X1  g695(.A1(new_n894_), .A2(new_n708_), .A3(new_n533_), .A4(new_n896_), .ZN(new_n897_));
  NOR4_X1   g696(.A1(new_n834_), .A2(new_n740_), .A3(new_n531_), .A4(new_n880_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n276_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT126), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n901_), .B(new_n897_), .C1(new_n898_), .C2(new_n276_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n834_), .A2(new_n531_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n321_), .A2(new_n511_), .A3(new_n444_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n737_), .A3(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G197gat), .ZN(G1352gat));
  AND3_X1   g706(.A1(new_n894_), .A2(new_n708_), .A3(new_n905_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G204gat), .B1(new_n909_), .B2(new_n650_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n644_), .A3(new_n390_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1353gat));
  XOR2_X1   g711(.A(KEYINPUT63), .B(G211gat), .Z(new_n913_));
  NAND4_X1  g712(.A1(new_n908_), .A2(KEYINPUT127), .A3(new_n565_), .A4(new_n913_), .ZN(new_n914_));
  OR2_X1    g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n908_), .B2(new_n565_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n904_), .A2(new_n565_), .A3(new_n905_), .A4(new_n913_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n914_), .B1(new_n916_), .B2(new_n919_), .ZN(G1354gat));
  AOI21_X1  g719(.A(G218gat), .B1(new_n908_), .B2(new_n614_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n680_), .A2(G218gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n908_), .B2(new_n922_), .ZN(G1355gat));
endmodule


