//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  OR2_X1    g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT9), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT10), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n202_), .B1(new_n211_), .B2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n223_), .A2(KEYINPUT9), .B1(new_n207_), .B2(new_n209_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n225_));
  AND2_X1   g024(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n225_), .B1(new_n228_), .B2(new_n215_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(new_n229_), .A3(KEYINPUT66), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n220_), .A2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n207_), .A2(new_n209_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n223_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n210_), .A2(new_n235_), .A3(new_n234_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT8), .A3(new_n223_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n244_));
  XOR2_X1   g043(.A(G71gat), .B(G78gat), .Z(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n246_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n231_), .A2(new_n242_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n246_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n249_), .B2(new_n247_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n240_), .A2(KEYINPUT8), .A3(new_n223_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT8), .B1(new_n240_), .B2(new_n223_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n220_), .A2(new_n230_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT12), .B1(new_n252_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n211_), .A2(new_n219_), .A3(new_n202_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT66), .B1(new_n224_), .B2(new_n229_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n239_), .B(new_n241_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT12), .B1(new_n266_), .B2(new_n251_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n260_), .A2(new_n263_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n251_), .B1(new_n231_), .B2(new_n242_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n257_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n263_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n267_), .B1(new_n274_), .B2(KEYINPUT12), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT67), .A3(new_n263_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G120gat), .B(G148gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n286_));
  INV_X1    g085(.A(new_n284_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n271_), .A2(new_n278_), .A3(new_n276_), .A4(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n279_), .A2(KEYINPUT69), .A3(new_n284_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT13), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT24), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  MUX2_X1   g095(.A(new_n295_), .B(KEYINPUT24), .S(new_n296_), .Z(new_n297_));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT23), .ZN(new_n299_));
  INV_X1    g098(.A(G190gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT26), .B1(new_n300_), .B2(KEYINPUT79), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G183gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G190gat), .ZN(new_n306_));
  OAI221_X1 g105(.A(new_n301_), .B1(new_n303_), .B2(new_n304_), .C1(KEYINPUT79), .C2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n304_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n302_), .A2(G183gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n297_), .B(new_n299_), .C1(new_n307_), .C2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n299_), .B1(G183gat), .B2(G190gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT80), .B(G176gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT22), .B(G169gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n294_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT81), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n311_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G71gat), .B(G99gat), .ZN(new_n322_));
  INV_X1    g121(.A(G43gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n321_), .A2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G227gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(G15gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT30), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n325_), .A2(new_n326_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT82), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT31), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n332_), .A2(new_n334_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(KEYINPUT82), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n343_), .B2(new_n335_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT89), .B(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G197gat), .ZN(new_n352_));
  INV_X1    g151(.A(G197gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT90), .B1(new_n353_), .B2(G204gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n350_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n353_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G197gat), .A2(G204gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT21), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n355_), .A2(KEYINPUT21), .A3(new_n356_), .A4(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n318_), .A2(new_n320_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT20), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n309_), .A2(new_n303_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n300_), .A2(KEYINPUT26), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n306_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n297_), .B(new_n299_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n316_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n367_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n366_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT93), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT93), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n380_), .A3(new_n377_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n368_), .A2(new_n373_), .A3(KEYINPUT95), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT95), .B1(new_n368_), .B2(new_n373_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n377_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n384_), .A2(KEYINPUT20), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n320_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n319_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT94), .B(new_n368_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT94), .B1(new_n321_), .B2(new_n368_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n383_), .B(new_n386_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n349_), .B1(new_n382_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n380_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n394_));
  AOI211_X1 g193(.A(KEYINPUT93), .B(new_n385_), .C1(new_n366_), .C2(new_n374_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n392_), .B(new_n349_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT83), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n400_), .A2(KEYINPUT3), .ZN(new_n401_));
  INV_X1    g200(.A(G141gat), .ZN(new_n402_));
  INV_X1    g201(.A(G148gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT2), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(G141gat), .A3(G148gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n404_), .A2(new_n406_), .B1(KEYINPUT84), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n400_), .A2(new_n409_), .A3(KEYINPUT3), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n401_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n401_), .A2(new_n408_), .A3(KEYINPUT85), .A4(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(KEYINPUT1), .B2(new_n416_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n416_), .A2(KEYINPUT1), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n402_), .A2(new_n403_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n399_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n420_), .A2(new_n421_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n419_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT86), .B1(new_n430_), .B2(new_n426_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n338_), .A3(new_n431_), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n430_), .A2(new_n338_), .A3(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT4), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n428_), .A2(new_n431_), .A3(new_n437_), .A4(new_n338_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G1gat), .B(G29gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G85gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT33), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n445_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n432_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n398_), .A2(new_n448_), .A3(new_n450_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n439_), .A2(new_n440_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n452_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n446_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n368_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n389_), .ZN(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT98), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n385_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n375_), .A2(new_n377_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT99), .B(new_n460_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n382_), .A2(new_n392_), .A3(new_n459_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n460_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT99), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n458_), .A2(new_n470_), .A3(new_n471_), .A4(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G22gat), .B(G50gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n428_), .A2(new_n431_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT29), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT87), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n483_));
  AOI211_X1 g282(.A(new_n483_), .B(KEYINPUT29), .C1(new_n428_), .C2(new_n431_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n479_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n421_), .B1(new_n420_), .B2(new_n427_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n430_), .A2(KEYINPUT86), .A3(new_n426_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n481_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n483_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(KEYINPUT87), .A3(new_n481_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n478_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G228gat), .A2(G233gat), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n368_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT29), .B1(new_n430_), .B2(new_n426_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n368_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(G228gat), .A3(G233gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G78gat), .B(G106gat), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n494_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n492_), .A2(KEYINPUT92), .A3(new_n500_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n492_), .A2(KEYINPUT92), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n502_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n485_), .A2(new_n491_), .A3(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n455_), .A2(new_n475_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n445_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n447_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n503_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT27), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n396_), .A2(KEYINPUT100), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT100), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n382_), .A2(new_n516_), .A3(new_n349_), .A4(new_n392_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n349_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n515_), .A2(new_n517_), .A3(KEYINPUT27), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n514_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n512_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n345_), .B1(new_n509_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT101), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT101), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n525_), .B(new_n345_), .C1(new_n509_), .C2(new_n522_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n344_), .A2(new_n511_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n521_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n508_), .A2(new_n503_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G8gat), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT75), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(G22gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n328_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G15gat), .A2(G22gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G1gat), .A2(G8gat), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n539_), .A2(new_n540_), .B1(KEYINPUT14), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n537_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G29gat), .B(G36gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n543_), .A2(new_n546_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n534_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n544_), .B(new_n545_), .Z(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n537_), .B(new_n542_), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n543_), .A2(new_n546_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(new_n533_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G169gat), .B(G197gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT77), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n549_), .A2(new_n556_), .A3(new_n563_), .A4(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n557_), .A2(KEYINPUT76), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT76), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n549_), .A2(new_n556_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n561_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n532_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n293_), .B1(new_n571_), .B2(KEYINPUT102), .ZN(new_n572_));
  INV_X1    g371(.A(new_n570_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n530_), .B1(new_n523_), .B2(KEYINPUT101), .ZN(new_n574_));
  AOI211_X1 g373(.A(KEYINPUT102), .B(new_n573_), .C1(new_n574_), .C2(new_n526_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n231_), .A2(new_n242_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n546_), .B(new_n551_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT71), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n580_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n266_), .B2(new_n550_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT72), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT71), .B1(new_n582_), .B2(new_n583_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n588_), .A2(KEYINPUT72), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n581_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OR3_X1    g392(.A1(new_n584_), .A2(new_n588_), .A3(new_n581_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT73), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT74), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n595_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n593_), .A2(new_n601_), .A3(new_n600_), .A4(new_n594_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT37), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(KEYINPUT37), .A3(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n251_), .B(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(new_n543_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n543_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n615_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(KEYINPUT17), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n615_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n610_), .A2(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n572_), .A2(new_n576_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(G1gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n458_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n605_), .A2(new_n606_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n293_), .A2(new_n573_), .ZN(new_n633_));
  AND4_X1   g432(.A1(new_n631_), .A2(new_n532_), .A3(new_n632_), .A4(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n511_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n628_), .A2(new_n629_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n636_), .A3(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n634_), .A2(new_n521_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G8gat), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n528_), .A2(G8gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n626_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n639_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n641_), .B(KEYINPUT39), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(KEYINPUT40), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1325gat));
  AOI21_X1  g449(.A(new_n328_), .B1(new_n634_), .B2(new_n344_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT41), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n626_), .A2(new_n328_), .A3(new_n344_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(new_n529_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n538_), .B1(new_n634_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT42), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n626_), .A2(new_n538_), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1327gat));
  AOI21_X1  g458(.A(new_n573_), .B1(new_n574_), .B2(new_n526_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n292_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n575_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n632_), .A2(new_n631_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n665_), .A2(G29gat), .A3(new_n511_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n633_), .A2(new_n624_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n605_), .A2(KEYINPUT37), .A3(new_n606_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n607_), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT43), .B(new_n670_), .C1(new_n574_), .C2(new_n526_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n532_), .B2(new_n610_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n668_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n532_), .A2(new_n610_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT43), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n532_), .A2(new_n672_), .A3(new_n610_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n667_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n458_), .B(new_n674_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n680_), .B2(G29gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n666_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  OAI211_X1 g483(.A(new_n521_), .B(new_n674_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n528_), .A2(G36gat), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n572_), .A2(new_n576_), .A3(new_n664_), .A4(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT45), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n663_), .A2(new_n690_), .A3(new_n664_), .A4(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n686_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n692_), .A3(KEYINPUT46), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n572_), .A2(new_n576_), .A3(new_n344_), .A4(new_n664_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(G43gat), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n674_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n344_), .A2(G43gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g503(.A(G50gat), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n701_), .A2(new_n705_), .A3(new_n529_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n665_), .B2(new_n529_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1331gat));
  INV_X1    g507(.A(new_n632_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n574_), .B2(new_n526_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n292_), .A2(new_n624_), .A3(new_n570_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n511_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n292_), .A2(new_n570_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n532_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n625_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n511_), .A2(G57gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1332gat));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719_));
  INV_X1    g518(.A(new_n712_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n521_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n721_), .B2(G64gat), .ZN(new_n722_));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT48), .B(new_n723_), .C1(new_n720_), .C2(new_n521_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n521_), .A2(new_n723_), .ZN(new_n725_));
  OAI22_X1  g524(.A1(new_n722_), .A2(new_n724_), .B1(new_n716_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT106), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n712_), .B2(new_n345_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n345_), .A2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n716_), .B2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n712_), .B2(new_n529_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n529_), .A2(G78gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n716_), .B2(new_n734_), .ZN(G1335gat));
  NAND3_X1  g534(.A1(new_n715_), .A2(new_n458_), .A3(new_n664_), .ZN(new_n736_));
  INV_X1    g535(.A(G85gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT107), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT107), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n676_), .A2(new_n677_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n292_), .A2(new_n631_), .A3(new_n570_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT108), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n458_), .A2(G85gat), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n739_), .A2(new_n740_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI221_X1 g547(.A(KEYINPUT109), .B1(new_n744_), .B2(new_n745_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1336gat));
  AND2_X1   g549(.A1(new_n715_), .A2(new_n664_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G92gat), .B1(new_n751_), .B2(new_n521_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n744_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n521_), .A2(G92gat), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT110), .Z(new_n755_));
  AOI21_X1  g554(.A(new_n752_), .B1(new_n753_), .B2(new_n755_), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n744_), .B2(new_n345_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n751_), .A2(new_n228_), .A3(new_n344_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n751_), .A2(new_n215_), .A3(new_n655_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n743_), .B(new_n655_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G106gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n761_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1339gat));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  NOR4_X1   g570(.A1(new_n655_), .A2(new_n521_), .A3(new_n345_), .A4(new_n511_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n260_), .A2(new_n268_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n275_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT12), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n774_), .B(new_n275_), .C1(new_n778_), .C2(new_n267_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n776_), .A2(new_n780_), .B1(new_n781_), .B2(new_n269_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT67), .B1(new_n277_), .B2(new_n263_), .ZN(new_n783_));
  NOR4_X1   g582(.A1(new_n778_), .A2(new_n270_), .A3(new_n267_), .A4(new_n275_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n284_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n284_), .A2(KEYINPUT56), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR4_X1   g592(.A1(new_n778_), .A2(new_n781_), .A3(new_n267_), .A4(new_n275_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT113), .B1(new_n277_), .B2(new_n263_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n779_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n271_), .A2(new_n781_), .A3(new_n278_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n789_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT114), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n788_), .A2(new_n793_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n533_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n554_), .A2(new_n555_), .A3(new_n534_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n561_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n565_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(new_n288_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT58), .B1(new_n800_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n773_), .B1(new_n807_), .B2(new_n670_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n287_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n809_));
  OAI22_X1  g608(.A1(KEYINPUT114), .A2(new_n798_), .B1(new_n809_), .B2(KEYINPUT56), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n791_), .A2(new_n792_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(KEYINPUT115), .A3(new_n610_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n806_), .B(KEYINPUT58), .C1(new_n810_), .C2(new_n811_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n808_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n791_), .B1(KEYINPUT56), .B2(new_n809_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n570_), .A2(new_n288_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n291_), .A2(new_n805_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n822_), .B2(new_n709_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n820_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n289_), .A2(new_n290_), .A3(new_n805_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT57), .B(new_n632_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n823_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n631_), .B1(new_n817_), .B2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n570_), .A2(new_n624_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n610_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n292_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(new_n292_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT59), .B(new_n772_), .C1(new_n828_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n834_), .A2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n823_), .A2(new_n826_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n816_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n670_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(KEYINPUT115), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n840_), .B1(new_n808_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n839_), .B1(new_n844_), .B2(new_n631_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT59), .B1(new_n845_), .B2(new_n772_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n771_), .B1(new_n838_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n772_), .B1(new_n828_), .B2(new_n836_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(KEYINPUT116), .A3(new_n837_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n573_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n848_), .B2(new_n573_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(KEYINPUT117), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1340gat));
  INV_X1    g659(.A(new_n848_), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n292_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n861_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n862_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n292_), .B1(new_n850_), .B2(new_n837_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n862_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n861_), .B2(new_n631_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n847_), .A2(new_n851_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(G127gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n631_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT120), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n869_), .B1(new_n870_), .B2(new_n873_), .ZN(G1342gat));
  INV_X1    g673(.A(G134gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n848_), .B2(new_n632_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT121), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n610_), .A2(G134gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n870_), .B2(new_n878_), .ZN(G1343gat));
  NOR2_X1   g678(.A1(new_n828_), .A2(new_n836_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n655_), .A2(new_n345_), .A3(new_n458_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n880_), .A2(new_n521_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n570_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n293_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT122), .B(G148gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1345gat));
  INV_X1    g686(.A(new_n882_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n888_), .B2(new_n624_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n882_), .A2(new_n890_), .A3(new_n631_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n889_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1346gat));
  INV_X1    g694(.A(G162gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n882_), .A2(new_n896_), .A3(new_n709_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n882_), .A2(new_n610_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n899_), .B2(new_n896_), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n880_), .A2(new_n528_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n527_), .A2(new_n529_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n570_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(G169gat), .B1(new_n903_), .B2(new_n573_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n314_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n906_), .B(new_n909_), .C1(new_n910_), .C2(new_n905_), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n901_), .A2(new_n293_), .A3(new_n902_), .ZN(new_n912_));
  INV_X1    g711(.A(G176gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  OR3_X1    g713(.A1(new_n912_), .A2(KEYINPUT125), .A3(new_n913_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n313_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n912_), .A2(KEYINPUT124), .A3(new_n313_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n914_), .A2(new_n915_), .B1(new_n918_), .B2(new_n919_), .ZN(G1349gat));
  NOR2_X1   g719(.A1(new_n903_), .A2(new_n624_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(G183gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n369_), .B2(new_n921_), .ZN(G1350gat));
  OR3_X1    g722(.A1(new_n903_), .A2(new_n632_), .A3(new_n371_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n904_), .A2(new_n610_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT126), .B1(new_n925_), .B2(G190gat), .ZN(new_n926_));
  OAI211_X1 g725(.A(KEYINPUT126), .B(G190gat), .C1(new_n903_), .C2(new_n670_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n924_), .B1(new_n926_), .B2(new_n928_), .ZN(G1351gat));
  NOR2_X1   g728(.A1(new_n512_), .A2(new_n344_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n901_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n573_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n353_), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n292_), .ZN(new_n934_));
  MUX2_X1   g733(.A(G204gat), .B(new_n351_), .S(new_n934_), .Z(G1353gat));
  AOI21_X1  g734(.A(new_n624_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT127), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n901_), .A2(new_n930_), .A3(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n938_), .B(new_n939_), .Z(G1354gat));
  OAI21_X1  g739(.A(G218gat), .B1(new_n931_), .B2(new_n670_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n632_), .A2(G218gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n931_), .B2(new_n942_), .ZN(G1355gat));
endmodule


