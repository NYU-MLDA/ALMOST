//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n207_), .B(new_n208_), .Z(new_n209_));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT87), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n210_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n211_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n213_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT88), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT2), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT3), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n214_), .A2(new_n218_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n219_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n213_), .B1(new_n216_), .B2(KEYINPUT1), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n212_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n225_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n209_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT4), .ZN(new_n231_));
  INV_X1    g030(.A(new_n229_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n207_), .B(new_n208_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n214_), .A2(new_n218_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n222_), .A2(new_n220_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(KEYINPUT4), .A3(new_n230_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT94), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n237_), .A2(new_n230_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(new_n241_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n206_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT33), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT95), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n241_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n231_), .A2(new_n238_), .A3(KEYINPUT95), .A4(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n205_), .B1(new_n243_), .B2(new_n241_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n249_), .B1(new_n231_), .B2(new_n238_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n243_), .A2(new_n241_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n205_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT33), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n246_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT19), .Z(new_n261_));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n262_));
  NOR2_X1   g061(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G169gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(G183gat), .A3(G190gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n264_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT83), .Z(new_n273_));
  INV_X1    g072(.A(KEYINPUT24), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(G169gat), .B2(G176gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT82), .B1(new_n278_), .B2(G183gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT25), .B(G183gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n277_), .B(new_n279_), .C1(new_n280_), .C2(KEYINPUT82), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n272_), .B(KEYINPUT83), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n274_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n268_), .A2(KEYINPUT84), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n268_), .A2(KEYINPUT84), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n266_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n271_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G197gat), .B(G204gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n290_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  OR3_X1    g093(.A1(new_n289_), .A2(new_n293_), .A3(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n262_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n269_), .B1(new_n274_), .B2(new_n272_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n275_), .A2(KEYINPUT90), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n275_), .A2(KEYINPUT90), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n273_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n277_), .A2(new_n280_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n264_), .B1(new_n287_), .B2(new_n270_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT91), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(KEYINPUT91), .B(new_n264_), .C1(new_n287_), .C2(new_n270_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n261_), .B(new_n297_), .C1(new_n309_), .C2(new_n296_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n296_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n309_), .B2(new_n296_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n312_), .B2(new_n261_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G8gat), .B(G36gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n318_), .B(new_n310_), .C1(new_n312_), .C2(new_n261_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n313_), .A2(KEYINPUT93), .A3(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n254_), .A2(new_n255_), .A3(new_n205_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n245_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n296_), .A2(KEYINPUT89), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n294_), .A2(new_n330_), .A3(new_n295_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n303_), .A2(new_n329_), .A3(new_n304_), .A4(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n261_), .B1(new_n297_), .B2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n312_), .B2(new_n261_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(KEYINPUT32), .ZN(new_n335_));
  MUX2_X1   g134(.A(new_n334_), .B(new_n313_), .S(new_n335_), .Z(new_n336_));
  AOI22_X1  g135(.A1(new_n259_), .A2(new_n325_), .B1(new_n328_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n288_), .B(KEYINPUT86), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G227gat), .A2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(G15gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT30), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n209_), .A2(KEYINPUT31), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n233_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G43gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .A4(new_n351_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n344_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n354_), .A3(new_n344_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n339_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n357_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n338_), .B1(new_n359_), .B2(new_n355_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n223_), .A2(new_n229_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n364_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n362_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n362_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n365_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n329_), .A2(new_n331_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n374_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n296_), .A2(new_n374_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n329_), .A2(new_n331_), .ZN(new_n384_));
  OAI211_X1 g183(.A(G228gat), .B(G233gat), .C1(new_n384_), .C2(new_n375_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n380_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n373_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n381_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n385_), .A2(new_n386_), .A3(new_n383_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n372_), .A4(new_n369_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n361_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n323_), .A2(new_n395_), .A3(new_n324_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n322_), .B(KEYINPUT27), .C1(new_n334_), .C2(new_n318_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n388_), .A2(new_n392_), .A3(new_n361_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n361_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n327_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n337_), .A2(new_n394_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G229gat), .A2(G233gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT15), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G29gat), .B(G36gat), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT71), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(KEYINPUT71), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G43gat), .B(G50gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n405_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(KEYINPUT15), .A3(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT76), .B(G15gat), .ZN(new_n417_));
  INV_X1    g216(.A(G22gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(G1gat), .ZN(new_n420_));
  INV_X1    g219(.A(G8gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT14), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G1gat), .B(G8gat), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n424_), .A3(new_n422_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n416_), .A2(KEYINPUT80), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n411_), .A2(new_n412_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n413_), .A2(new_n415_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(new_n430_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n404_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n431_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n428_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n432_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n403_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT81), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G113gat), .B(G141gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G169gat), .B(G197gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n442_), .A2(KEYINPUT81), .A3(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n402_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT96), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT13), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G120gat), .B(G148gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT5), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G176gat), .B(G204gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(G230gat), .A2(G233gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT64), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT64), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G85gat), .ZN(new_n471_));
  INV_X1    g270(.A(G92gat), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n471_), .A2(new_n472_), .A3(KEYINPUT9), .ZN(new_n473_));
  XOR2_X1   g272(.A(G85gat), .B(G92gat), .Z(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(KEYINPUT9), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT10), .B(G99gat), .Z(new_n476_));
  INV_X1    g275(.A(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n470_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n466_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n484_), .B(new_n485_), .C1(G99gat), .C2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n487_), .B(new_n477_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n474_), .B1(new_n483_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT8), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n486_), .A2(new_n488_), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT8), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n474_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n480_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G57gat), .B(G64gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT11), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT66), .B(G71gat), .ZN(new_n501_));
  INV_X1    g300(.A(G78gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n501_), .B(G78gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n499_), .A2(KEYINPUT11), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n498_), .A2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n460_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT12), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n498_), .B2(new_n508_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n460_), .B1(new_n498_), .B2(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n479_), .A2(KEYINPUT68), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT68), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n470_), .A2(new_n475_), .A3(new_n517_), .A4(new_n478_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n474_), .ZN(new_n520_));
  AOI211_X1 g319(.A(KEYINPUT8), .B(new_n520_), .C1(new_n470_), .C2(new_n494_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n496_), .B1(new_n495_), .B2(new_n474_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT67), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n493_), .A2(new_n524_), .A3(new_n497_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n519_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n508_), .A2(new_n513_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n514_), .B(new_n515_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n459_), .B1(new_n512_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n512_), .A2(new_n528_), .A3(new_n459_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT69), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n531_), .B2(KEYINPUT69), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n530_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n534_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n454_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(KEYINPUT13), .A3(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G190gat), .B(G218gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT36), .Z(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n498_), .B2(new_n431_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n549_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT35), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n551_), .B(new_n555_), .C1(new_n526_), .C2(new_n435_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n550_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n479_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n559_), .B1(new_n560_), .B2(new_n438_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n519_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT67), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n524_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n561_), .B1(new_n565_), .B2(new_n416_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(new_n555_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n547_), .B1(new_n558_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n416_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(new_n557_), .A3(new_n555_), .A4(new_n551_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n556_), .A2(KEYINPUT72), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n551_), .B1(new_n526_), .B2(new_n435_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n554_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n573_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n574_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n568_), .B(new_n569_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n557_), .B1(new_n566_), .B2(new_n555_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n556_), .A2(KEYINPUT72), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n577_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT73), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n573_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT74), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT75), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n568_), .A2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT75), .B(new_n547_), .C1(new_n558_), .C2(new_n567_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n583_), .A2(new_n589_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n581_), .B1(new_n593_), .B2(KEYINPUT37), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n428_), .B(new_n595_), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n508_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G127gat), .B(G155gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n597_), .A2(KEYINPUT17), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n604_));
  AND4_X1   g403(.A1(new_n604_), .A2(new_n597_), .A3(KEYINPUT17), .A4(new_n602_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n597_), .A2(new_n604_), .B1(KEYINPUT17), .B2(new_n602_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT79), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n594_), .A2(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n453_), .A2(new_n543_), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n420_), .A3(new_n328_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n587_), .A2(new_n588_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n568_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n402_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(new_n607_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n542_), .A2(new_n450_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n327_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n612_), .A2(new_n613_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n621_), .A3(new_n622_), .ZN(G1324gat));
  NAND3_X1  g422(.A1(new_n611_), .A2(new_n421_), .A3(new_n398_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n398_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G8gat), .B1(new_n620_), .B2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g429(.A(new_n620_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n361_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n341_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT41), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n611_), .A2(new_n341_), .A3(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT97), .ZN(G1326gat));
  NOR2_X1   g436(.A1(new_n389_), .A2(new_n393_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G22gat), .B1(new_n620_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT98), .Z(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT42), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n611_), .A2(new_n418_), .A3(new_n638_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(KEYINPUT42), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(G1327gat));
  INV_X1    g444(.A(new_n616_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n609_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n542_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n453_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n328_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n609_), .A2(new_n539_), .A3(new_n451_), .A4(new_n541_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n593_), .A2(KEYINPUT37), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n402_), .A3(new_n580_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n594_), .A2(new_n657_), .A3(new_n402_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n653_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n652_), .B1(new_n659_), .B2(KEYINPUT99), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n661_), .B(new_n653_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n651_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n653_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n658_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n657_), .B1(new_n594_), .B2(new_n402_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n661_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n665_), .B(KEYINPUT99), .C1(new_n666_), .C2(new_n667_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(KEYINPUT100), .A3(new_n652_), .A4(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n664_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n659_), .A2(KEYINPUT44), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n328_), .A2(G29gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n650_), .B1(new_n676_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n453_), .A2(new_n679_), .A3(new_n398_), .A4(new_n648_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT45), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n674_), .A2(new_n398_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n663_), .B2(new_n671_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(new_n679_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n684_), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT46), .B1(new_n684_), .B2(KEYINPUT101), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  NAND2_X1  g486(.A1(new_n663_), .A2(new_n671_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(G43gat), .A3(new_n632_), .A4(new_n674_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G43gat), .B1(new_n649_), .B2(new_n632_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT47), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n689_), .A2(new_n694_), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1330gat));
  INV_X1    g495(.A(G50gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n638_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT102), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n649_), .A2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n673_), .A2(new_n639_), .A3(new_n675_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n697_), .ZN(G1331gat));
  NOR2_X1   g501(.A1(new_n543_), .A2(new_n451_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n402_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n704_), .A2(new_n594_), .A3(new_n609_), .ZN(new_n705_));
  INV_X1    g504(.A(G57gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n328_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n607_), .B(KEYINPUT79), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n708_), .A3(new_n617_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT103), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(new_n328_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n711_), .B2(new_n706_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n710_), .B2(new_n398_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT48), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n705_), .A2(new_n713_), .A3(new_n398_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n710_), .B2(new_n632_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT49), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n705_), .A2(new_n718_), .A3(new_n632_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1334gat));
  AOI21_X1  g521(.A(new_n502_), .B1(new_n710_), .B2(new_n638_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT50), .Z(new_n724_));
  NAND2_X1  g523(.A1(new_n638_), .A2(new_n502_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT104), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n705_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n704_), .A2(new_n647_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n471_), .A3(new_n328_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n609_), .B(new_n703_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n327_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1336gat));
  NAND3_X1  g532(.A1(new_n729_), .A2(new_n472_), .A3(new_n398_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G92gat), .B1(new_n731_), .B2(new_n625_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1337gat));
  NAND3_X1  g535(.A1(new_n729_), .A2(new_n632_), .A3(new_n476_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT105), .Z(new_n738_));
  OAI21_X1  g537(.A(G99gat), .B1(new_n731_), .B2(new_n361_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n731_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n477_), .B1(new_n744_), .B2(new_n638_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n746_));
  INV_X1    g545(.A(new_n647_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n639_), .A2(G106gat), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n703_), .A2(new_n747_), .A3(new_n402_), .A4(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT106), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n746_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n752_), .A2(KEYINPUT108), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755_));
  INV_X1    g554(.A(new_n753_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n750_), .B1(new_n745_), .B2(KEYINPUT52), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n743_), .B1(new_n754_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT108), .B1(new_n752_), .B2(new_n753_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n757_), .A3(new_n755_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n742_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n646_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n429_), .A2(new_n432_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT80), .B1(new_n416_), .B2(new_n428_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n436_), .A2(KEYINPUT112), .A3(new_n432_), .A4(new_n429_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n403_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n440_), .A2(new_n404_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n447_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n446_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n773_), .B(new_n774_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n448_), .A2(new_n449_), .A3(new_n531_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n526_), .A2(new_n527_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(KEYINPUT55), .A3(new_n514_), .A4(new_n515_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n514_), .B(new_n509_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n460_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n528_), .A2(new_n781_), .ZN(new_n782_));
  AND4_X1   g581(.A1(KEYINPUT110), .A2(new_n778_), .A3(new_n780_), .A4(new_n782_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n528_), .A2(new_n781_), .B1(new_n779_), .B2(new_n460_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n784_), .B2(new_n778_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n458_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n782_), .B(new_n780_), .C1(new_n789_), .C2(new_n528_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n784_), .A2(KEYINPUT110), .A3(new_n778_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n458_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n776_), .B1(new_n788_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n775_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n448_), .A2(new_n449_), .A3(new_n531_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n458_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n787_), .B(new_n459_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(KEYINPUT111), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n765_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n773_), .A2(new_n531_), .A3(new_n774_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n773_), .A2(KEYINPUT113), .A3(new_n531_), .A4(new_n774_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(KEYINPUT114), .A2(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI221_X1 g611(.A(new_n809_), .B1(KEYINPUT114), .B2(KEYINPUT58), .C1(new_n800_), .C2(new_n801_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n594_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n773_), .A2(new_n774_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n540_), .B2(new_n536_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n802_), .B2(KEYINPUT111), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n796_), .A2(new_n797_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n646_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n804_), .B(new_n814_), .C1(new_n819_), .C2(KEYINPUT57), .ZN(new_n820_));
  INV_X1    g619(.A(new_n607_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n610_), .A2(new_n450_), .A3(new_n543_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT54), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n610_), .A2(new_n824_), .A3(new_n450_), .A4(new_n543_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n820_), .A2(new_n821_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n625_), .A2(new_n328_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n400_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n451_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n609_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n823_), .A2(new_n825_), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT59), .B(new_n830_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT115), .B1(new_n831_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(KEYINPUT59), .C1(new_n826_), .C2(new_n830_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n450_), .B(new_n836_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n833_), .B1(new_n841_), .B2(new_n832_), .ZN(G1340gat));
  XNOR2_X1  g641(.A(KEYINPUT116), .B(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n543_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n831_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n843_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n543_), .B(new_n836_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g646(.A(G127gat), .B1(new_n831_), .B2(new_n708_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n836_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT117), .B(G127gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n821_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n848_), .B1(new_n849_), .B2(new_n851_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n831_), .A2(new_n853_), .A3(new_n646_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n594_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n855_), .B(new_n836_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n856_), .B2(new_n853_), .ZN(G1343gat));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  INV_X1    g657(.A(new_n399_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n827_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n826_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n804_), .A2(new_n814_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n616_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n764_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n607_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n823_), .A2(new_n825_), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT118), .B(new_n860_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n451_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n542_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g672(.A1(new_n869_), .A2(new_n708_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877_));
  AOI21_X1  g676(.A(G162gat), .B1(new_n869_), .B2(new_n646_), .ZN(new_n878_));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n855_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n862_), .B2(new_n868_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n877_), .B1(new_n878_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n869_), .A2(new_n880_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n616_), .B1(new_n862_), .B2(new_n868_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n884_), .B(KEYINPUT119), .C1(G162gat), .C2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n886_), .ZN(G1347gat));
  NAND2_X1  g686(.A1(new_n834_), .A2(new_n835_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n625_), .A2(new_n328_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n828_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT120), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT22), .B(G169gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n451_), .A2(new_n894_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT121), .Z(new_n896_));
  NAND3_X1  g695(.A1(new_n888_), .A2(new_n451_), .A3(new_n891_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(new_n898_), .A3(G169gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(G169gat), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n893_), .A2(new_n896_), .B1(new_n899_), .B2(new_n900_), .ZN(G1348gat));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n892_), .B(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n542_), .ZN(new_n904_));
  INV_X1    g703(.A(G176gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n826_), .A2(new_n638_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n543_), .A2(new_n890_), .A3(new_n905_), .A4(new_n361_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n904_), .A2(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n609_), .A2(new_n890_), .A3(new_n361_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G183gat), .B1(new_n906_), .B2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n821_), .A2(new_n280_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n903_), .B2(new_n911_), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n893_), .B2(new_n855_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n903_), .A2(new_n277_), .A3(new_n646_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1351gat));
  NOR3_X1   g714(.A1(new_n826_), .A2(new_n859_), .A3(new_n890_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916_), .B2(new_n451_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n917_), .A2(KEYINPUT123), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(KEYINPUT123), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(G197gat), .A3(new_n451_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n916_), .A2(KEYINPUT122), .A3(G197gat), .A4(new_n451_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n918_), .A2(new_n919_), .B1(new_n922_), .B2(new_n923_), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n916_), .A2(new_n542_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n607_), .A2(new_n927_), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT124), .Z(new_n929_));
  NAND2_X1  g728(.A1(new_n916_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n931_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT126), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n933_), .B(new_n935_), .ZN(G1354gat));
  AND3_X1   g735(.A1(new_n916_), .A2(G218gat), .A3(new_n594_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n916_), .A2(new_n646_), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n938_), .A2(KEYINPUT127), .ZN(new_n939_));
  AOI21_X1  g738(.A(G218gat), .B1(new_n938_), .B2(KEYINPUT127), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n937_), .B1(new_n939_), .B2(new_n940_), .ZN(G1355gat));
endmodule


