//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n202_), .B(new_n203_), .C1(new_n209_), .C2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n218_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(KEYINPUT65), .ZN(new_n220_));
  OAI21_X1  g019(.A(G85gat), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n214_), .B1(new_n202_), .B2(KEYINPUT9), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n225_), .B2(new_n206_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n224_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n221_), .B(new_n222_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n215_), .A2(new_n216_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n217_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n230_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n217_), .A2(new_n237_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT12), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT12), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n230_), .A2(new_n242_), .A3(new_n238_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G230gat), .A2(G233gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(new_n240_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n245_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G120gat), .B(G148gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G176gat), .B(G204gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n253_), .B(new_n254_), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n246_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT13), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n257_), .B(new_n258_), .C1(KEYINPUT68), .C2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G229gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G29gat), .B(G36gat), .ZN(new_n266_));
  INV_X1    g065(.A(G43gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(G50gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G22gat), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G8gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n269_), .B(KEYINPUT15), .ZN(new_n278_));
  INV_X1    g077(.A(new_n276_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n265_), .B(new_n277_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n269_), .A2(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n265_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G113gat), .B(G141gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G197gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT70), .ZN(new_n287_));
  INV_X1    g086(.A(G169gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n280_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n264_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n279_), .B(new_n237_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G231gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT17), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT16), .B(G183gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G211gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n299_), .A2(new_n300_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(KEYINPUT17), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT22), .B(G169gat), .ZN(new_n309_));
  INV_X1    g108(.A(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n317_), .A3(KEYINPUT73), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n319_), .A3(KEYINPUT23), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n318_), .B(new_n320_), .C1(G183gat), .C2(G190gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT96), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n322_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n313_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT95), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n315_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT75), .B1(new_n314_), .B2(KEYINPUT23), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n331_), .A2(new_n316_), .A3(G183gat), .A4(G190gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n314_), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n288_), .A2(new_n310_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n335_), .A2(KEYINPUT24), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT94), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT94), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(new_n339_), .A3(new_n336_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n312_), .A2(KEYINPUT24), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT93), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT26), .B(G190gat), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT25), .B(G183gat), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n344_), .A2(new_n335_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n327_), .B1(new_n341_), .B2(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n334_), .A2(new_n339_), .A3(new_n336_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n339_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n348_), .B(new_n327_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n326_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT97), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT21), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT87), .ZN(new_n360_));
  OR2_X1    g159(.A1(G211gat), .A2(G218gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G211gat), .A2(G218gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n358_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n356_), .A2(new_n357_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n365_), .B(new_n368_), .C1(new_n366_), .C2(new_n358_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n354_), .A2(new_n355_), .A3(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n348_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT95), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n325_), .B1(new_n376_), .B2(new_n352_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT97), .B1(new_n377_), .B2(new_n372_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT88), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n372_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n370_), .A2(KEYINPUT88), .A3(new_n371_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G183gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT71), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT71), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(G183gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n387_), .A3(KEYINPUT25), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n345_), .A2(KEYINPUT72), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n391_));
  INV_X1    g190(.A(G190gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(KEYINPUT26), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n335_), .A2(KEYINPUT24), .A3(new_n312_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n318_), .A2(new_n320_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .A4(new_n336_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n385_), .A2(new_n387_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n334_), .B1(G190gat), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n313_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n379_), .B1(new_n383_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n374_), .A2(new_n378_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT92), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT19), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n382_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT88), .B1(new_n370_), .B2(new_n371_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n379_), .B1(new_n412_), .B2(new_n402_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n377_), .B2(new_n372_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT18), .B(G64gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G92gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n409_), .A2(new_n420_), .A3(new_n415_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT78), .B(G113gat), .ZN(new_n424_));
  INV_X1    g223(.A(G120gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n424_), .A2(new_n425_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428_));
  OR3_X1    g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432_));
  INV_X1    g231(.A(G141gat), .ZN(new_n433_));
  INV_X1    g232(.A(G148gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G155gat), .A2(G162gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT81), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT1), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n435_), .B(new_n436_), .C1(new_n438_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n435_), .B1(new_n442_), .B2(KEYINPUT3), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT2), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n436_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(new_n433_), .A3(new_n434_), .A4(KEYINPUT82), .ZN(new_n447_));
  NAND3_X1  g246(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n443_), .A2(new_n445_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n439_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n441_), .B1(new_n450_), .B2(new_n438_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n431_), .A2(new_n432_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n431_), .B(new_n451_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n452_), .B(new_n454_), .C1(new_n455_), .C2(new_n432_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n431_), .B(new_n451_), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n453_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT0), .B(G57gat), .ZN(new_n459_));
  INV_X1    g258(.A(G85gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G1gat), .B(G29gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT33), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n456_), .A2(new_n458_), .A3(new_n467_), .A4(new_n464_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n452_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n457_), .B2(KEYINPUT4), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n464_), .B1(new_n470_), .B2(new_n453_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n457_), .A2(new_n454_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n466_), .A2(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n422_), .A2(new_n423_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT98), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n456_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n464_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT99), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  AND4_X1   g279(.A1(new_n479_), .A2(new_n456_), .A3(new_n458_), .A4(new_n464_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n326_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n413_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n408_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n420_), .A2(KEYINPUT32), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n482_), .B(new_n488_), .C1(new_n416_), .C2(new_n487_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n422_), .A2(KEYINPUT98), .A3(new_n473_), .A4(new_n423_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n476_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n431_), .B(KEYINPUT31), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n397_), .A2(new_n495_), .A3(new_n401_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n402_), .A2(KEYINPUT30), .ZN(new_n499_));
  INV_X1    g298(.A(new_n494_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n397_), .A2(new_n495_), .A3(new_n401_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G15gat), .B(G43gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G227gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G71gat), .B(G99gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  AND3_X1   g306(.A1(new_n498_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT79), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n511_));
  INV_X1    g310(.A(new_n507_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n496_), .A2(new_n497_), .A3(new_n494_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n500_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n498_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n511_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n493_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT79), .B1(new_n508_), .B2(new_n509_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n493_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n492_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n515_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n520_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n515_), .A2(new_n516_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n493_), .B1(new_n525_), .B2(KEYINPUT79), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n524_), .A2(new_n526_), .A3(KEYINPUT80), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n522_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n529_));
  INV_X1    g328(.A(G233gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT84), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(G228gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(G228gat), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT85), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n451_), .A2(KEYINPUT29), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n381_), .A2(new_n535_), .A3(new_n536_), .A4(new_n382_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n535_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(new_n372_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G78gat), .B(G106gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT89), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n545_), .A3(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G22gat), .B(G50gat), .ZN(new_n548_));
  OR3_X1    g347(.A1(new_n451_), .A2(KEYINPUT29), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n451_), .B2(KEYINPUT29), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n529_), .B1(new_n547_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n542_), .B2(new_n541_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n546_), .A2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n546_), .A2(new_n558_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n547_), .A2(new_n529_), .A3(new_n554_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n491_), .A2(new_n528_), .A3(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n562_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(new_n555_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n518_), .A2(new_n521_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n561_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT27), .ZN(new_n572_));
  INV_X1    g371(.A(new_n423_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n420_), .B1(new_n409_), .B2(new_n415_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n482_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n486_), .A2(new_n421_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(KEYINPUT27), .A3(new_n423_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n579_), .ZN(new_n580_));
  AOI211_X1 g379(.A(new_n295_), .B(new_n308_), .C1(new_n565_), .C2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n230_), .A2(new_n269_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n217_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n586_));
  OAI221_X1 g385(.A(new_n583_), .B1(KEYINPUT35), .B2(new_n585_), .C1(new_n278_), .C2(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(KEYINPUT35), .B(new_n585_), .C1(new_n582_), .C2(KEYINPUT69), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G134gat), .ZN(new_n593_));
  INV_X1    g392(.A(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n589_), .A2(new_n590_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n595_), .B(KEYINPUT36), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n600_), .A3(new_n590_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT37), .B1(new_n603_), .B2(new_n596_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n581_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT101), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n607_), .B(KEYINPUT100), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n610_), .A2(new_n613_), .A3(new_n271_), .A4(new_n482_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n603_), .A2(new_n596_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n581_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n576_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n615_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n619_), .A3(new_n620_), .ZN(G1324gat));
  NAND2_X1  g420(.A1(new_n575_), .A2(new_n578_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n610_), .A2(new_n613_), .A3(new_n272_), .A4(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n618_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT102), .B(G8gat), .C1(new_n618_), .C2(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(KEYINPUT103), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT103), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n630_), .A2(KEYINPUT103), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n627_), .A2(new_n632_), .A3(new_n633_), .A4(new_n628_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n623_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n623_), .A2(KEYINPUT40), .A3(new_n631_), .A4(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  NOR3_X1   g438(.A1(new_n611_), .A2(G15gat), .A3(new_n528_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G15gat), .B1(new_n618_), .B2(new_n528_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT41), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1326gat));
  OAI21_X1  g442(.A(G22gat), .B1(new_n618_), .B2(new_n564_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT42), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n564_), .A2(G22gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT104), .Z(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n611_), .B2(new_n647_), .ZN(G1327gat));
  AOI21_X1  g447(.A(new_n617_), .B1(new_n565_), .B2(new_n580_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n308_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n295_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n482_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n565_), .A2(new_n580_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n605_), .ZN(new_n656_));
  AOI211_X1 g455(.A(KEYINPUT43), .B(new_n606_), .C1(new_n565_), .C2(new_n580_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n651_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT44), .B(new_n651_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(G29gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n653_), .B1(new_n663_), .B2(new_n482_), .ZN(G1328gat));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n665_), .A2(KEYINPUT107), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(new_n622_), .A3(new_n661_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G36gat), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n667_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n652_), .A2(new_n673_), .A3(new_n622_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n676_), .A2(new_n677_), .B1(KEYINPUT107), .B2(new_n665_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n666_), .B1(new_n672_), .B2(new_n678_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n667_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT105), .B1(new_n667_), .B2(G36gat), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n666_), .B(new_n678_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n679_), .A2(new_n683_), .ZN(G1329gat));
  INV_X1    g483(.A(new_n528_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n652_), .A2(new_n267_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n662_), .A2(new_n569_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(G43gat), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g489(.A(G50gat), .B1(new_n652_), .B2(new_n563_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n563_), .A2(G50gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n662_), .B2(new_n692_), .ZN(G1331gat));
  AOI211_X1 g492(.A(new_n294_), .B(new_n264_), .C1(new_n565_), .C2(new_n580_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n602_), .A2(new_n604_), .A3(new_n650_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT108), .Z(new_n698_));
  AOI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n482_), .ZN(new_n699_));
  OR2_X1    g498(.A1(KEYINPUT109), .A2(G57gat), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n694_), .A2(new_n617_), .A3(new_n650_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n576_), .B2(KEYINPUT109), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n699_), .B1(new_n700_), .B2(new_n703_), .ZN(G1332gat));
  OR3_X1    g503(.A1(new_n697_), .A2(G64gat), .A3(new_n624_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n622_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G64gat), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT48), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT48), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n705_), .B1(new_n710_), .B2(new_n711_), .ZN(G1333gat));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n701_), .B2(new_n685_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT49), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n697_), .A2(G71gat), .A3(new_n528_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1334gat));
  INV_X1    g516(.A(G78gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n701_), .B2(new_n563_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT50), .Z(new_n720_));
  NAND2_X1  g519(.A1(new_n563_), .A2(new_n718_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT111), .Z(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n697_), .B2(new_n722_), .ZN(G1335gat));
  NOR3_X1   g522(.A1(new_n264_), .A2(new_n650_), .A3(new_n294_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n649_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n482_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n656_), .A2(new_n657_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n724_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n576_), .A2(new_n460_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1336gat));
  AOI21_X1  g531(.A(G92gat), .B1(new_n726_), .B2(new_n622_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT65), .B(G92gat), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n624_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n730_), .B2(new_n735_), .ZN(G1337gat));
  OAI21_X1  g535(.A(G99gat), .B1(new_n729_), .B2(new_n528_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n726_), .A2(new_n225_), .A3(new_n569_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n563_), .B(new_n724_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n743_), .B2(new_n206_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n726_), .A2(new_n206_), .A3(new_n563_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n746_), .A2(new_n751_), .A3(new_n748_), .A4(new_n749_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1339gat));
  OAI21_X1  g554(.A(G113gat), .B1(new_n293_), .B2(KEYINPUT120), .ZN(new_n756_));
  OR2_X1    g555(.A1(KEYINPUT120), .A2(G113gat), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n622_), .A2(new_n576_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n570_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n244_), .A2(new_n245_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n246_), .A2(KEYINPUT55), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n244_), .A2(new_n766_), .A3(new_n245_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n768_), .B2(new_n255_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT55), .B(new_n248_), .C1(new_n241_), .C2(new_n243_), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n770_), .A2(new_n771_), .B1(new_n245_), .B2(new_n244_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n256_), .A3(new_n762_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n769_), .A2(new_n294_), .A3(new_n258_), .A4(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n256_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n293_), .B1(new_n777_), .B2(new_n763_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n778_), .A2(KEYINPUT116), .A3(new_n258_), .A4(new_n773_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n283_), .B(new_n277_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n289_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n282_), .A2(new_n265_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n783_), .A2(KEYINPUT117), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT117), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n259_), .A2(new_n784_), .A3(new_n290_), .A4(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n776_), .A2(new_n779_), .A3(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n787_), .A2(KEYINPUT57), .A3(new_n617_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT57), .B1(new_n787_), .B2(new_n617_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n777_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n256_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(KEYINPUT118), .A3(new_n793_), .ZN(new_n794_));
  AND4_X1   g593(.A1(new_n290_), .A2(new_n784_), .A3(new_n258_), .A4(new_n785_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n796_), .A3(new_n791_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n794_), .A2(KEYINPUT58), .A3(new_n795_), .A4(new_n797_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n605_), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n650_), .B1(new_n790_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n264_), .A2(new_n293_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n696_), .B2(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n695_), .A2(KEYINPUT54), .A3(new_n805_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT59), .B(new_n761_), .C1(new_n803_), .C2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n787_), .A2(new_n617_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n787_), .A2(KEYINPUT57), .A3(new_n617_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n802_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n809_), .B1(new_n816_), .B2(new_n308_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n811_), .B1(new_n817_), .B2(new_n760_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n810_), .A2(new_n818_), .A3(KEYINPUT119), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT119), .B1(new_n810_), .B2(new_n818_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n756_), .B(new_n757_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n817_), .A2(new_n293_), .A3(new_n760_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n822_), .A2(G113gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT121), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n821_), .A2(new_n826_), .A3(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1340gat));
  NAND2_X1  g627(.A1(new_n810_), .A2(new_n818_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n264_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n831_), .A2(KEYINPUT122), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(KEYINPUT122), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(G120gat), .A3(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n817_), .A2(new_n760_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n425_), .B1(new_n264_), .B2(KEYINPUT60), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n835_), .B(new_n836_), .C1(KEYINPUT60), .C2(new_n425_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n835_), .B2(new_n650_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n819_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n820_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n308_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n839_), .B1(new_n842_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g642(.A(new_n617_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G134gat), .B1(new_n835_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n606_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g646(.A1(new_n817_), .A2(new_n566_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n758_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n293_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT123), .B(G141gat), .Z(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1344gat));
  NOR2_X1   g651(.A1(new_n849_), .A2(new_n264_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n434_), .ZN(G1345gat));
  NOR2_X1   g653(.A1(new_n849_), .A2(new_n308_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT61), .B(G155gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  NOR3_X1   g656(.A1(new_n849_), .A2(new_n594_), .A3(new_n606_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n848_), .A2(new_n844_), .A3(new_n758_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n594_), .B2(new_n859_), .ZN(G1347gat));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n817_), .A2(new_n563_), .A3(new_n624_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n528_), .A2(new_n482_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n294_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n861_), .B1(new_n866_), .B2(G169gat), .ZN(new_n867_));
  AOI211_X1 g666(.A(KEYINPUT62), .B(new_n288_), .C1(new_n865_), .C2(new_n294_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n294_), .A2(new_n309_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT124), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n867_), .A2(new_n868_), .B1(new_n864_), .B2(new_n870_), .ZN(G1348gat));
  NOR2_X1   g670(.A1(new_n864_), .A2(new_n264_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n310_), .ZN(G1349gat));
  NOR2_X1   g672(.A1(new_n864_), .A2(new_n308_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n347_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n876_), .B(new_n877_), .C1(new_n398_), .C2(new_n874_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n877_), .B2(new_n876_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n864_), .B2(new_n606_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n844_), .A2(new_n346_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n864_), .B2(new_n881_), .ZN(G1351gat));
  NOR2_X1   g681(.A1(new_n624_), .A2(new_n482_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n848_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n293_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT126), .B(G197gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1352gat));
  INV_X1    g686(.A(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n830_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g689(.A1(new_n884_), .A2(new_n308_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n891_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT63), .B(G211gat), .Z(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(new_n893_), .ZN(G1354gat));
  NAND3_X1  g693(.A1(new_n888_), .A2(KEYINPUT127), .A3(new_n844_), .ZN(new_n895_));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n884_), .B2(new_n617_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n896_), .A3(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n888_), .A2(G218gat), .A3(new_n605_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1355gat));
endmodule


