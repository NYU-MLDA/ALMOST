//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n989_,
    new_n990_, new_n991_, new_n993_, new_n994_, new_n996_, new_n997_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1013_, new_n1014_, new_n1015_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  OR3_X1    g008(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT83), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n211_), .B1(new_n213_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT26), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT26), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n222_), .B(new_n224_), .C1(new_n225_), .C2(G183gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n228_));
  OAI21_X1  g027(.A(G183gat), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT81), .B(G183gat), .C1(new_n227_), .C2(new_n228_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n226_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n220_), .B1(new_n233_), .B2(KEYINPUT82), .ZN(new_n234_));
  INV_X1    g033(.A(new_n226_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT80), .B(KEYINPUT25), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT81), .B1(new_n236_), .B2(G183gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n232_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n218_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n212_), .A2(new_n218_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT85), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n208_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT22), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n206_), .B1(new_n251_), .B2(G169gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT84), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(G169gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(KEYINPUT84), .A3(G169gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n250_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n258_));
  OAI22_X1  g057(.A1(new_n234_), .A2(new_n241_), .B1(new_n249_), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G211gat), .B(G218gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT93), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n260_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n264_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n262_), .A2(new_n263_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT92), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n265_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  AOI211_X1 g071(.A(new_n202_), .B(new_n204_), .C1(new_n259_), .C2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n208_), .B(KEYINPUT101), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n254_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT23), .B1(new_n214_), .B2(new_n216_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n213_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI221_X1 g078(.A(new_n274_), .B1(G176gat), .B2(new_n276_), .C1(new_n279_), .C2(new_n243_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT100), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT98), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n223_), .A2(G190gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n221_), .A2(KEYINPUT26), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT25), .B(G183gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT98), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT99), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n209_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n210_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n242_), .A2(new_n292_), .A3(new_n245_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(new_n289_), .B2(new_n209_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n282_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n289_), .A2(new_n209_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT99), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n298_), .A2(KEYINPUT100), .A3(new_n291_), .A4(new_n293_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n281_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n272_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n273_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n259_), .B2(new_n272_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n280_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n306_), .B2(new_n272_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n204_), .B(KEYINPUT97), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n303_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G8gat), .B(G36gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n303_), .B(new_n317_), .C1(new_n307_), .C2(new_n309_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(KEYINPUT103), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT103), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n310_), .A2(new_n321_), .A3(new_n315_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT91), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n272_), .B2(KEYINPUT94), .ZN(new_n327_));
  INV_X1    g126(.A(G155gat), .ZN(new_n328_));
  INV_X1    g127(.A(G162gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AND3_X1   g129(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT89), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT89), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n330_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n344_), .A2(new_n347_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n334_), .A2(new_n341_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n345_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(new_n342_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n339_), .A2(KEYINPUT1), .B1(new_n328_), .B2(new_n329_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n337_), .A2(new_n356_), .A3(new_n338_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n351_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n272_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n327_), .A2(new_n361_), .ZN(new_n362_));
  OAI221_X1 g161(.A(new_n272_), .B1(KEYINPUT94), .B2(new_n326_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(KEYINPUT95), .A3(new_n368_), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n364_), .A2(KEYINPUT95), .A3(new_n365_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n359_), .A2(new_n372_), .A3(new_n360_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n357_), .A3(new_n330_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n353_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n334_), .A2(new_n341_), .A3(new_n350_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT28), .B1(new_n378_), .B2(KEYINPUT29), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n380_), .A2(new_n382_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n371_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(KEYINPUT90), .A3(new_n383_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n369_), .A2(new_n370_), .A3(new_n386_), .A4(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n366_), .A2(KEYINPUT96), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n364_), .A2(new_n391_), .A3(new_n365_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n384_), .A2(new_n385_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .A4(new_n368_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n301_), .B1(new_n305_), .B2(new_n280_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n396_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n204_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n280_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT107), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n280_), .B(KEYINPUT107), .C1(new_n294_), .C2(new_n295_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n301_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n202_), .B1(new_n259_), .B2(new_n272_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n398_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n315_), .B1(new_n397_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(KEYINPUT27), .A3(new_n318_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n323_), .A2(new_n395_), .A3(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G127gat), .B(G134gat), .Z(new_n409_));
  XOR2_X1   g208(.A(G113gat), .B(G120gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n209_), .B(new_n210_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n233_), .A2(KEYINPUT82), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n254_), .A2(new_n253_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n256_), .A3(new_n206_), .A4(new_n275_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n208_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n242_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n243_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n244_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n417_), .B1(new_n420_), .B2(KEYINPUT85), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n413_), .A2(new_n414_), .B1(new_n421_), .B2(new_n248_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT30), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(G15gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G43gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G99gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n422_), .A2(KEYINPUT30), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n423_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n430_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT87), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT31), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n423_), .A2(new_n431_), .A3(new_n432_), .A4(new_n434_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n411_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT31), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n409_), .B(new_n410_), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G1gat), .B(G29gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT105), .B(KEYINPUT0), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n378_), .A2(new_n454_), .A3(new_n444_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G225gat), .A2(G233gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n444_), .B1(new_n351_), .B2(new_n358_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n376_), .A2(new_n377_), .A3(new_n411_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT104), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT104), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n378_), .A2(new_n462_), .A3(new_n444_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n458_), .B1(new_n464_), .B2(KEYINPUT4), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n457_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n453_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n456_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n454_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n468_), .B(new_n452_), .C1(new_n469_), .C2(new_n458_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n408_), .A2(new_n447_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n469_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n455_), .A2(new_n456_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n452_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n461_), .A2(KEYINPUT106), .A3(new_n463_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT106), .B1(new_n461_), .B2(new_n463_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n457_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(KEYINPUT33), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n470_), .A2(KEYINPUT33), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(new_n319_), .B2(new_n322_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n303_), .B(new_n485_), .C1(new_n307_), .C2(new_n309_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n471_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n307_), .A2(new_n309_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n405_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n485_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT108), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n202_), .B1(new_n422_), .B2(new_n301_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n301_), .B2(new_n300_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n493_), .A2(new_n308_), .B1(new_n302_), .B2(new_n273_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n494_), .A2(new_n485_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT108), .ZN(new_n496_));
  INV_X1    g295(.A(new_n485_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n397_), .B2(new_n405_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n491_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n395_), .B1(new_n484_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n471_), .B1(new_n389_), .B2(new_n394_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n323_), .A2(new_n502_), .A3(new_n407_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n472_), .B1(new_n504_), .B2(new_n447_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G29gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT75), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n509_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n509_), .B(KEYINPUT15), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n518_), .B(new_n519_), .C1(new_n521_), .C2(new_n517_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n509_), .B(new_n517_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n519_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n525_), .A2(KEYINPUT78), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(KEYINPUT78), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n522_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G113gat), .B(G141gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT79), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n522_), .B(new_n532_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n505_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G64gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G57gat), .ZN(new_n540_));
  INV_X1    g339(.A(G57gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(G64gat), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n540_), .A2(new_n542_), .A3(KEYINPUT69), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT69), .B1(new_n540_), .B2(new_n542_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT11), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n541_), .A2(G64gat), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n539_), .A2(G57gat), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT11), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n540_), .A2(new_n542_), .A3(KEYINPUT69), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G71gat), .B(G78gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT11), .B(new_n553_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(G106gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT6), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT6), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(G99gat), .A3(G106gat), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n560_), .A2(new_n561_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT9), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT65), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT65), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT9), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n568_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT66), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OAI211_X1 g380(.A(KEYINPUT67), .B(new_n566_), .C1(new_n576_), .C2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n563_), .A2(new_n565_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n584_));
  OR3_X1    g383(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT8), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n575_), .A2(KEYINPUT68), .A3(new_n567_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n582_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n576_), .A2(new_n581_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT67), .B1(new_n592_), .B2(new_n566_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n557_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n555_), .A2(new_n556_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(new_n588_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT8), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT67), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n576_), .A2(new_n581_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n566_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n595_), .A2(new_n599_), .A3(new_n603_), .A4(new_n582_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n594_), .A2(KEYINPUT12), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n557_), .B(new_n606_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT64), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT70), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n594_), .A2(new_n604_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n610_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(KEYINPUT70), .A3(new_n611_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G120gat), .B(G148gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n614_), .A2(new_n616_), .A3(new_n617_), .A4(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT72), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT70), .B1(new_n608_), .B2(new_n611_), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n613_), .B(new_n610_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n628_), .A2(KEYINPUT72), .A3(new_n616_), .A4(new_n622_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n616_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n622_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n630_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n595_), .B(new_n517_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT17), .ZN(new_n643_));
  XOR2_X1   g442(.A(G127gat), .B(G155gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT16), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n642_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(KEYINPUT17), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT37), .ZN(new_n652_));
  INV_X1    g451(.A(new_n591_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n603_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n520_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n509_), .A3(new_n603_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(G232gat), .A2(G233gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT34), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(KEYINPUT35), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(KEYINPUT35), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT74), .Z(new_n661_));
  INV_X1    g460(.A(KEYINPUT76), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n655_), .A2(new_n656_), .A3(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n661_), .A2(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n655_), .A2(new_n667_), .A3(new_n656_), .A4(new_n663_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G190gat), .B(G218gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(G134gat), .B(G162gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT36), .Z(new_n672_));
  NAND4_X1  g471(.A1(new_n666_), .A2(KEYINPUT77), .A3(new_n668_), .A4(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n666_), .A2(new_n668_), .A3(new_n672_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT77), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n671_), .A2(KEYINPUT36), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n652_), .B(new_n673_), .C1(new_n676_), .C2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n674_), .A2(KEYINPUT37), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(new_n679_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n638_), .A2(new_n651_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n538_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n471_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n685_), .A2(G1gat), .A3(new_n686_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT38), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT38), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n389_), .A2(new_n394_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n496_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n691_));
  AND4_X1   g490(.A1(new_n496_), .A2(new_n498_), .A3(new_n471_), .A4(new_n486_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n482_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n694_), .A2(new_n480_), .B1(new_n478_), .B2(new_n475_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n318_), .A2(KEYINPUT103), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n494_), .A2(new_n317_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n322_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n690_), .B1(new_n693_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n503_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n447_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n447_), .A2(new_n471_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n323_), .A2(new_n407_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(new_n395_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n673_), .B1(new_n676_), .B2(new_n679_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT109), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(new_n673_), .C1(new_n676_), .C2(new_n679_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n651_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n536_), .B(new_n715_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n708_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G1gat), .B1(new_n718_), .B2(new_n686_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n688_), .A2(new_n689_), .A3(new_n719_), .ZN(G1324gat));
  INV_X1    g519(.A(KEYINPUT40), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT39), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n722_), .B(G8gat), .C1(new_n718_), .C2(new_n706_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n505_), .A2(new_n713_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n705_), .A3(new_n717_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n727_), .A2(KEYINPUT111), .A3(new_n722_), .A4(G8gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G8gat), .B1(new_n718_), .B2(new_n706_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT39), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n730_), .B2(KEYINPUT39), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n729_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n685_), .A2(G8gat), .A3(new_n706_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n721_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n735_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n732_), .A2(new_n733_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT40), .B(new_n737_), .C1(new_n738_), .C2(new_n729_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1325gat));
  NOR3_X1   g539(.A1(new_n685_), .A2(G15gat), .A3(new_n447_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT112), .Z(new_n742_));
  INV_X1    g541(.A(new_n718_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n447_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n425_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n747_), .A3(new_n748_), .ZN(G1326gat));
  OAI21_X1  g548(.A(G22gat), .B1(new_n718_), .B2(new_n395_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT42), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n395_), .A2(G22gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n685_), .B2(new_n752_), .ZN(G1327gat));
  NOR3_X1   g552(.A1(new_n714_), .A2(new_n638_), .A3(new_n715_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n538_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(G29gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n471_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n536_), .B(new_n651_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n680_), .A2(new_n682_), .A3(KEYINPUT114), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT114), .B1(new_n680_), .B2(new_n682_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n762_), .B1(new_n708_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n683_), .A2(new_n762_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n505_), .A2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT44), .B(new_n761_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT115), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n744_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n765_), .B1(new_n771_), .B2(new_n472_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT43), .ZN(new_n773_));
  INV_X1    g572(.A(new_n767_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n708_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(KEYINPUT44), .A4(new_n761_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n770_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n761_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n686_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI211_X1 g581(.A(KEYINPUT116), .B(new_n757_), .C1(new_n779_), .C2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n759_), .B(KEYINPUT113), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n777_), .B1(new_n786_), .B2(KEYINPUT44), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n772_), .A2(KEYINPUT43), .B1(new_n708_), .B2(new_n774_), .ZN(new_n788_));
  NOR4_X1   g587(.A1(new_n788_), .A2(new_n785_), .A3(KEYINPUT115), .A4(new_n781_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n782_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(new_n790_), .B2(G29gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n758_), .B1(new_n783_), .B2(new_n791_), .ZN(G1328gat));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n793_));
  INV_X1    g592(.A(G36gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n706_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n779_), .B2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n705_), .A2(KEYINPUT117), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n705_), .A2(KEYINPUT117), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n794_), .ZN(new_n800_));
  OR3_X1    g599(.A1(new_n755_), .A2(KEYINPUT45), .A3(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT45), .B1(new_n755_), .B2(new_n800_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n793_), .B1(new_n796_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n705_), .B1(new_n786_), .B2(KEYINPUT44), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n770_), .B2(new_n778_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT46), .B(new_n803_), .C1(new_n807_), .C2(new_n794_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(G1329gat));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n755_), .A2(new_n447_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n787_), .A2(new_n789_), .ZN(new_n812_));
  OAI211_X1 g611(.A(G43gat), .B(new_n744_), .C1(new_n786_), .C2(KEYINPUT44), .ZN(new_n813_));
  OAI221_X1 g612(.A(new_n810_), .B1(G43gat), .B2(new_n811_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n770_), .B2(new_n778_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n811_), .A2(G43gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT47), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(G1330gat));
  OR3_X1    g617(.A1(new_n755_), .A2(G50gat), .A3(new_n395_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n395_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n779_), .A2(KEYINPUT118), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G50gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT118), .B1(new_n779_), .B2(new_n820_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(G1331gat));
  NOR2_X1   g623(.A1(new_n505_), .A2(new_n536_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n683_), .A2(new_n651_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n638_), .A3(new_n826_), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT119), .Z(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n541_), .A3(new_n471_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n726_), .A2(new_n537_), .A3(new_n638_), .A4(new_n715_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G57gat), .B1(new_n830_), .B2(new_n686_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1332gat));
  INV_X1    g631(.A(new_n799_), .ZN(new_n833_));
  OAI21_X1  g632(.A(G64gat), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT48), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n799_), .A2(new_n539_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT120), .Z(new_n837_));
  NAND2_X1  g636(.A1(new_n828_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(G1333gat));
  INV_X1    g638(.A(G71gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n828_), .A2(new_n840_), .A3(new_n744_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G71gat), .B1(new_n830_), .B2(new_n447_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT49), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1334gat));
  INV_X1    g643(.A(G78gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n828_), .A2(new_n845_), .A3(new_n690_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G78gat), .B1(new_n830_), .B2(new_n395_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT50), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1335gat));
  NAND2_X1  g648(.A1(new_n638_), .A2(new_n651_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n714_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n825_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(G85gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n471_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n850_), .A2(new_n536_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n788_), .A2(new_n686_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n858_), .B2(new_n854_), .ZN(G1336gat));
  INV_X1    g658(.A(G92gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n853_), .A2(new_n860_), .A3(new_n705_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n788_), .A2(new_n833_), .A3(new_n857_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1337gat));
  NAND2_X1  g662(.A1(new_n744_), .A2(new_n560_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n852_), .A2(new_n864_), .B1(KEYINPUT121), .B2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n776_), .A2(new_n744_), .A3(new_n856_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(G99gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(KEYINPUT121), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n868_), .B(new_n869_), .Z(G1338gat));
  NAND3_X1  g669(.A1(new_n853_), .A2(new_n561_), .A3(new_n690_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n776_), .A2(new_n690_), .A3(new_n856_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n872_), .A2(new_n873_), .A3(G106gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n872_), .B2(G106gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n871_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT53), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n878_), .B(new_n871_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1339gat));
  NOR3_X1   g679(.A1(new_n408_), .A2(new_n447_), .A3(new_n686_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(KEYINPUT59), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n626_), .A2(new_n627_), .A3(KEYINPUT55), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n608_), .A2(KEYINPUT55), .A3(new_n611_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n611_), .B2(new_n608_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n632_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n887_), .A2(KEYINPUT56), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(KEYINPUT56), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n888_), .A2(new_n536_), .A3(new_n630_), .A4(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n532_), .B1(new_n523_), .B2(new_n519_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n521_), .A2(new_n517_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n518_), .A2(new_n524_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n535_), .A2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT122), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n630_), .A2(new_n633_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n713_), .B1(new_n890_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n896_), .A2(new_n888_), .A3(new_n630_), .A4(new_n889_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n889_), .A2(new_n630_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n905_), .A2(KEYINPUT58), .A3(new_n896_), .A4(new_n888_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n683_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n715_), .B1(new_n901_), .B2(new_n907_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n635_), .A2(new_n637_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n537_), .A3(new_n826_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n883_), .B1(new_n908_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n907_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n890_), .A2(new_n898_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n714_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n900_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n904_), .A2(KEYINPUT123), .A3(new_n683_), .A4(new_n906_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n899_), .A2(KEYINPUT57), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n915_), .A2(new_n918_), .A3(new_n919_), .A4(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n912_), .B1(new_n921_), .B2(new_n651_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n882_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n536_), .B(new_n913_), .C1(new_n923_), .C2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(G113gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n921_), .A2(new_n651_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n912_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n881_), .ZN(new_n930_));
  OR3_X1    g729(.A1(new_n930_), .A2(G113gat), .A3(new_n537_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n926_), .A2(new_n931_), .ZN(G1340gat));
  OAI211_X1 g731(.A(new_n638_), .B(new_n913_), .C1(new_n923_), .C2(new_n924_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G120gat), .ZN(new_n934_));
  INV_X1    g733(.A(G120gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n909_), .B2(KEYINPUT60), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n923_), .B(new_n936_), .C1(KEYINPUT60), .C2(new_n935_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(G1341gat));
  AOI21_X1  g737(.A(G127gat), .B1(new_n923_), .B2(new_n715_), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n908_), .A2(new_n912_), .ZN(new_n940_));
  AOI22_X1  g739(.A1(new_n930_), .A2(KEYINPUT59), .B1(new_n940_), .B2(new_n883_), .ZN(new_n941_));
  INV_X1    g740(.A(G127gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n715_), .B2(KEYINPUT124), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(KEYINPUT124), .B2(new_n942_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n939_), .B1(new_n941_), .B2(new_n944_), .ZN(G1342gat));
  OAI211_X1 g744(.A(new_n683_), .B(new_n913_), .C1(new_n923_), .C2(new_n924_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(G134gat), .ZN(new_n947_));
  OR3_X1    g746(.A1(new_n930_), .A2(G134gat), .A3(new_n714_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1343gat));
  NOR2_X1   g748(.A1(new_n922_), .A2(new_n744_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n799_), .A2(new_n686_), .A3(new_n395_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  OAI21_X1  g751(.A(G141gat), .B1(new_n952_), .B2(new_n537_), .ZN(new_n953_));
  INV_X1    g752(.A(G141gat), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n950_), .A2(new_n954_), .A3(new_n536_), .A4(new_n951_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1344gat));
  OAI21_X1  g755(.A(G148gat), .B1(new_n952_), .B2(new_n909_), .ZN(new_n957_));
  INV_X1    g756(.A(G148gat), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n950_), .A2(new_n958_), .A3(new_n638_), .A4(new_n951_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n959_), .ZN(G1345gat));
  XNOR2_X1  g759(.A(KEYINPUT61), .B(G155gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n952_), .B2(new_n651_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n961_), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n950_), .A2(new_n715_), .A3(new_n951_), .A4(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1346gat));
  INV_X1    g764(.A(new_n952_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n763_), .A2(new_n764_), .A3(new_n329_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n950_), .A2(new_n713_), .A3(new_n951_), .ZN(new_n968_));
  AOI22_X1  g767(.A1(new_n966_), .A2(new_n967_), .B1(new_n968_), .B2(new_n329_), .ZN(G1347gat));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n908_), .A2(new_n912_), .ZN(new_n971_));
  AND2_X1   g770(.A1(new_n799_), .A2(new_n704_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(new_n395_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n971_), .A2(new_n537_), .A3(new_n973_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n970_), .B1(new_n974_), .B2(new_n205_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n973_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n940_), .A2(new_n536_), .A3(new_n976_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n977_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n974_), .A2(new_n254_), .A3(new_n275_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n975_), .A2(new_n978_), .A3(new_n979_), .ZN(G1348gat));
  NOR2_X1   g779(.A1(new_n971_), .A2(new_n973_), .ZN(new_n981_));
  AOI21_X1  g780(.A(G176gat), .B1(new_n981_), .B2(new_n638_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n929_), .A2(KEYINPUT125), .A3(new_n395_), .ZN(new_n983_));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n984_), .B1(new_n922_), .B2(new_n690_), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n983_), .A2(new_n985_), .A3(new_n972_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n909_), .A2(new_n206_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n982_), .B1(new_n986_), .B2(new_n987_), .ZN(G1349gat));
  NAND4_X1  g787(.A1(new_n983_), .A2(new_n985_), .A3(new_n715_), .A4(new_n972_), .ZN(new_n989_));
  INV_X1    g788(.A(G183gat), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n651_), .A2(new_n287_), .ZN(new_n991_));
  AOI22_X1  g790(.A1(new_n989_), .A2(new_n990_), .B1(new_n981_), .B2(new_n991_), .ZN(G1350gat));
  NAND4_X1  g791(.A1(new_n981_), .A2(new_n286_), .A3(new_n288_), .A4(new_n713_), .ZN(new_n993_));
  AND2_X1   g792(.A1(new_n981_), .A2(new_n683_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n994_), .B2(new_n221_), .ZN(G1351gat));
  AND2_X1   g794(.A1(new_n799_), .A2(new_n502_), .ZN(new_n996_));
  NAND4_X1  g795(.A1(new_n929_), .A2(new_n447_), .A3(new_n536_), .A4(new_n996_), .ZN(new_n997_));
  XNOR2_X1  g796(.A(new_n997_), .B(G197gat), .ZN(G1352gat));
  XNOR2_X1  g797(.A(KEYINPUT126), .B(G204gat), .ZN(new_n999_));
  INV_X1    g798(.A(new_n999_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n950_), .A2(new_n996_), .ZN(new_n1001_));
  OAI21_X1  g800(.A(new_n1000_), .B1(new_n1001_), .B2(new_n909_), .ZN(new_n1002_));
  NAND4_X1  g801(.A1(new_n950_), .A2(new_n638_), .A3(new_n996_), .A4(new_n999_), .ZN(new_n1003_));
  NAND2_X1  g802(.A1(new_n1002_), .A2(new_n1003_), .ZN(G1353gat));
  NOR2_X1   g803(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1005_));
  XNOR2_X1  g804(.A(new_n1005_), .B(KEYINPUT127), .ZN(new_n1006_));
  INV_X1    g805(.A(new_n1006_), .ZN(new_n1007_));
  AOI21_X1  g806(.A(new_n651_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1008_));
  INV_X1    g807(.A(new_n1008_), .ZN(new_n1009_));
  OAI21_X1  g808(.A(new_n1007_), .B1(new_n1001_), .B2(new_n1009_), .ZN(new_n1010_));
  NAND4_X1  g809(.A1(new_n950_), .A2(new_n996_), .A3(new_n1006_), .A4(new_n1008_), .ZN(new_n1011_));
  NAND2_X1  g810(.A1(new_n1010_), .A2(new_n1011_), .ZN(G1354gat));
  AND3_X1   g811(.A1(new_n950_), .A2(new_n683_), .A3(new_n996_), .ZN(new_n1013_));
  INV_X1    g812(.A(G218gat), .ZN(new_n1014_));
  NAND2_X1  g813(.A1(new_n713_), .A2(new_n1014_), .ZN(new_n1015_));
  OAI22_X1  g814(.A1(new_n1013_), .A2(new_n1014_), .B1(new_n1001_), .B2(new_n1015_), .ZN(G1355gat));
endmodule


