//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT89), .Z(new_n212_));
  OAI211_X1 g011(.A(new_n202_), .B(new_n204_), .C1(new_n210_), .C2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n209_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n203_), .B(KEYINPUT3), .Z(new_n215_));
  XOR2_X1   g014(.A(new_n202_), .B(KEYINPUT2), .Z(new_n216_));
  OAI211_X1 g015(.A(new_n207_), .B(new_n214_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G127gat), .B(G134gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n220_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT86), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n221_), .A2(new_n223_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n218_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(KEYINPUT4), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n231_), .B1(new_n235_), .B2(new_n230_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G1gat), .B(G29gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G85gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n236_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT99), .ZN(new_n244_));
  OR3_X1    g043(.A1(new_n218_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT28), .B1(new_n218_), .B2(KEYINPUT29), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G22gat), .B(G50gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n218_), .A2(KEYINPUT29), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT91), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G197gat), .B(G204gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n250_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(G228gat), .A2(G233gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n259_), .B2(KEYINPUT90), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n250_), .B(new_n259_), .C1(KEYINPUT90), .C2(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(KEYINPUT93), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n265_), .A2(new_n268_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n249_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT94), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n249_), .B(KEYINPUT94), .C1(new_n269_), .C2(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n265_), .A2(KEYINPUT92), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n265_), .A2(KEYINPUT92), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n266_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n249_), .B1(new_n266_), .B2(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT82), .B(G176gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT83), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n284_), .A2(new_n285_), .B1(G169gat), .B2(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT84), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(KEYINPUT23), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(KEYINPUT23), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n289_), .B1(new_n290_), .B2(new_n287_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  OAI221_X1 g091(.A(new_n286_), .B1(new_n285_), .B2(new_n284_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT24), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n294_), .A2(KEYINPUT24), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT25), .B(G183gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  AOI211_X1 g098(.A(new_n295_), .B(new_n297_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n290_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(new_n301_), .A3(KEYINPUT30), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(KEYINPUT85), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(KEYINPUT85), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G71gat), .B(G99gat), .ZN(new_n311_));
  INV_X1    g110(.A(G43gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(G15gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n313_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n310_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n307_), .A2(new_n317_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n226_), .B(KEYINPUT31), .Z(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n316_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(new_n319_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(KEYINPUT87), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n321_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n324_), .A2(new_n319_), .A3(new_n323_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n281_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n273_), .A2(new_n274_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n328_), .A2(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n244_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT20), .B1(new_n302_), .B2(new_n259_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n336_), .A2(KEYINPUT95), .ZN(new_n337_));
  INV_X1    g136(.A(new_n291_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n300_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n284_), .A2(new_n296_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT96), .ZN(new_n341_));
  INV_X1    g140(.A(new_n290_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n292_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n340_), .A2(KEYINPUT96), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n339_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n259_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n336_), .B2(KEYINPUT95), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n337_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n302_), .A2(new_n259_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n349_), .B(KEYINPUT20), .C1(new_n259_), .C2(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  MUX2_X1   g151(.A(new_n348_), .B(new_n350_), .S(new_n352_), .Z(new_n353_));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT18), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n352_), .B1(new_n337_), .B2(new_n347_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n350_), .A2(new_n352_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n357_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT100), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT100), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT27), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n357_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n363_), .A2(KEYINPUT27), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n357_), .A2(KEYINPUT32), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n353_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n360_), .A2(new_n361_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n373_), .B(new_n243_), .C1(new_n374_), .C2(new_n372_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n236_), .A2(KEYINPUT33), .A3(new_n242_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT33), .B1(new_n236_), .B2(new_n242_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n241_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n235_), .B2(new_n230_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT97), .B1(new_n363_), .B2(new_n369_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n363_), .A2(KEYINPUT97), .A3(new_n369_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n375_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n330_), .A2(new_n326_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(new_n281_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n335_), .A2(new_n371_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G229gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(KEYINPUT77), .B(G8gat), .Z(new_n390_));
  INV_X1    g189(.A(G1gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT14), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT76), .B(G15gat), .ZN(new_n393_));
  INV_X1    g192(.A(G22gat), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G1gat), .B(G8gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n392_), .A2(new_n395_), .A3(new_n396_), .A4(new_n398_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G29gat), .B(G36gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G43gat), .B(G50gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n389_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407_));
  INV_X1    g206(.A(new_n402_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n405_), .B(KEYINPUT15), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT15), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n405_), .B(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n412_), .A2(new_n402_), .A3(KEYINPUT81), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n406_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n402_), .B(new_n405_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n389_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G141gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G169gat), .B(G197gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n387_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G64gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G57gat), .ZN(new_n426_));
  INV_X1    g225(.A(G57gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G64gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n428_), .A3(KEYINPUT11), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT68), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G57gat), .B(G64gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT11), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G71gat), .B(G78gat), .Z(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(KEYINPUT11), .B2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(new_n430_), .A3(new_n433_), .A4(new_n435_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(G85gat), .A2(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n445_));
  INV_X1    g244(.A(G99gat), .ZN(new_n446_));
  INV_X1    g245(.A(G106gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n448_), .B(new_n449_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT67), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n454_), .A2(new_n456_), .A3(new_n451_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n444_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n451_), .A2(new_n453_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n448_), .A2(new_n459_), .A3(new_n449_), .A4(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(KEYINPUT66), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n441_), .A2(new_n463_), .A3(new_n442_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n461_), .B2(KEYINPUT66), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n458_), .A2(KEYINPUT8), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT10), .B(G99gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT65), .B(G85gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT9), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G92gat), .ZN(new_n470_));
  OAI22_X1  g269(.A1(G106gat), .A2(new_n467_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n459_), .B(new_n460_), .C1(new_n443_), .C2(new_n469_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n440_), .B(KEYINPUT12), .C1(new_n466_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n437_), .A2(new_n439_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n473_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n462_), .A2(new_n465_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n451_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n448_), .A2(new_n449_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n450_), .A2(new_n451_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n463_), .B1(new_n483_), .B2(new_n444_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n475_), .B(new_n476_), .C1(new_n477_), .C2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n474_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT69), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G230gat), .A2(G233gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT64), .Z(new_n489_));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n457_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT8), .B1(new_n491_), .B2(new_n443_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n462_), .A2(new_n465_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n473_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n490_), .B1(new_n494_), .B2(new_n475_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n486_), .A2(new_n487_), .A3(new_n489_), .A4(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n489_), .A3(new_n485_), .A4(new_n474_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT69), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n500_));
  INV_X1    g299(.A(new_n489_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n485_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n494_), .A2(new_n475_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G120gat), .B(G148gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT5), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G176gat), .B(G204gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .A4(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n496_), .A2(new_n498_), .A3(new_n504_), .A4(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT70), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n499_), .A2(new_n504_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n508_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n513_), .B(new_n515_), .C1(KEYINPUT71), .C2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n515_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n517_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G190gat), .B(G218gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G134gat), .B(G162gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT34), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n476_), .B1(new_n477_), .B2(new_n484_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n405_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n494_), .A2(new_n412_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT35), .B(new_n528_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534_));
  INV_X1    g333(.A(new_n528_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n494_), .A2(new_n405_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n534_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n529_), .A2(new_n409_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n526_), .B1(new_n541_), .B2(KEYINPUT74), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT74), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n533_), .A2(new_n543_), .A3(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT37), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n524_), .A2(new_n525_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT72), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n533_), .A2(new_n540_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n526_), .B1(new_n533_), .B2(new_n540_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n551_), .A2(KEYINPUT73), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n551_), .B2(KEYINPUT73), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT37), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT75), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n550_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT78), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n402_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n440_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT80), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT17), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n564_), .B(new_n570_), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n563_), .A2(KEYINPUT17), .A3(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n559_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n424_), .A2(new_n521_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT101), .ZN(new_n577_));
  INV_X1    g376(.A(new_n521_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n575_), .ZN(new_n579_));
  NOR4_X1   g378(.A1(new_n387_), .A2(new_n423_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT101), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n391_), .A3(new_n244_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n583_), .A2(KEYINPUT38), .A3(new_n391_), .A4(new_n244_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n545_), .A2(new_n549_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n387_), .A2(new_n574_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n423_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n521_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n244_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n587_), .A3(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(new_n371_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n577_), .A2(new_n598_), .A3(new_n582_), .A4(new_n390_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n590_), .A2(new_n598_), .A3(new_n593_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n600_), .A2(new_n601_), .A3(G8gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n600_), .B2(G8gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(G1325gat));
  INV_X1    g405(.A(new_n385_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G15gat), .B1(new_n594_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT41), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n576_), .A2(G15gat), .A3(new_n607_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1326gat));
  NAND3_X1  g410(.A1(new_n580_), .A2(new_n394_), .A3(new_n281_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G22gat), .B1(new_n594_), .B2(new_n332_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT42), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT42), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(G1327gat));
  NOR2_X1   g415(.A1(new_n573_), .A2(new_n588_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n521_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n424_), .A2(new_n618_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n619_), .A2(G29gat), .A3(new_n595_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n592_), .A2(new_n573_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n556_), .A2(new_n558_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n387_), .A2(KEYINPUT43), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n334_), .B1(new_n385_), .B2(new_n332_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n371_), .A3(new_n595_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n384_), .A2(new_n386_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n625_), .B1(new_n629_), .B2(new_n559_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n622_), .B1(new_n624_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT43), .B1(new_n387_), .B2(new_n623_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(new_n625_), .A3(new_n559_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(KEYINPUT44), .A3(new_n622_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n621_), .B1(new_n638_), .B2(new_n244_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n633_), .A2(new_n621_), .A3(new_n244_), .A4(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G29gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n620_), .B1(new_n639_), .B2(new_n641_), .ZN(G1328gat));
  INV_X1    g441(.A(KEYINPUT46), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(KEYINPUT104), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n633_), .A2(new_n598_), .A3(new_n637_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G36gat), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n371_), .A2(G36gat), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n424_), .A2(new_n648_), .A3(new_n618_), .A4(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n629_), .A2(new_n591_), .A3(new_n618_), .A4(new_n649_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT45), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n643_), .A2(KEYINPUT104), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n645_), .B1(new_n647_), .B2(new_n656_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n644_), .B(new_n655_), .C1(new_n646_), .C2(G36gat), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1329gat));
  NAND4_X1  g458(.A1(new_n633_), .A2(G43gat), .A3(new_n333_), .A4(new_n637_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n312_), .B1(new_n619_), .B2(new_n607_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g462(.A(new_n619_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G50gat), .B1(new_n664_), .B2(new_n281_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n281_), .A2(G50gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n638_), .B2(new_n666_), .ZN(G1331gat));
  NAND2_X1  g466(.A1(new_n578_), .A2(new_n423_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n590_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(G57gat), .A3(new_n244_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT106), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n629_), .A2(new_n423_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(new_n521_), .A3(new_n579_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT105), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G57gat), .B1(new_n676_), .B2(new_n244_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n672_), .A2(new_n677_), .ZN(G1332gat));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n425_), .A3(new_n598_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n425_), .B1(new_n670_), .B2(new_n598_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT48), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(G1333gat));
  OR2_X1    g483(.A1(new_n607_), .A2(G71gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n590_), .A2(new_n385_), .A3(new_n669_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT49), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G71gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G71gat), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n675_), .A2(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  OAI221_X1 g491(.A(new_n692_), .B1(new_n688_), .B2(new_n689_), .C1(new_n675_), .C2(new_n685_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1334gat));
  INV_X1    g493(.A(G78gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n670_), .B2(new_n281_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT50), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n281_), .A2(new_n695_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT108), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n698_), .A2(new_n699_), .B1(new_n675_), .B2(new_n701_), .ZN(G1335gat));
  NAND2_X1  g501(.A1(new_n578_), .A2(new_n617_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n673_), .A2(KEYINPUT109), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT109), .B1(new_n673_), .B2(new_n703_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n244_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n636_), .A2(new_n574_), .A3(new_n669_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(new_n595_), .A3(new_n468_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1336gat));
  INV_X1    g509(.A(G92gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n711_), .A3(new_n598_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G92gat), .B1(new_n708_), .B2(new_n371_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1337gat));
  OAI21_X1  g513(.A(G99gat), .B1(new_n708_), .B2(new_n607_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n328_), .A2(new_n329_), .A3(new_n467_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n706_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n718_), .A2(KEYINPUT110), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(KEYINPUT110), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1338gat));
  XNOR2_X1  g521(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n669_), .A2(new_n574_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n332_), .B(new_n724_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT52), .B1(new_n725_), .B2(new_n447_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n636_), .A2(new_n281_), .A3(new_n574_), .A4(new_n669_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(G106gat), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n281_), .A2(new_n447_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n723_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n723_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n732_), .B(new_n735_), .C1(new_n726_), .C2(new_n729_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  INV_X1    g536(.A(KEYINPUT59), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n623_), .A2(new_n521_), .A3(new_n423_), .A4(new_n573_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(KEYINPUT112), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n575_), .A2(new_n423_), .A3(new_n521_), .A4(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n423_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n497_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n474_), .A2(new_n485_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT12), .B1(new_n529_), .B2(new_n440_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n501_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT113), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n501_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n749_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n496_), .A2(new_n498_), .A3(new_n748_), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n747_), .B(new_n509_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n753_), .A2(new_n755_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n749_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n757_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n508_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n746_), .B1(new_n758_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT114), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n746_), .B(new_n765_), .C1(new_n758_), .C2(new_n762_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n419_), .B1(new_n415_), .B2(new_n388_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n410_), .A2(new_n413_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n389_), .B1(new_n408_), .B2(new_n530_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT115), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n767_), .B(new_n772_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n420_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n518_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n764_), .A2(new_n766_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n588_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(KEYINPUT57), .A3(new_n588_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n774_), .B1(new_n512_), .B2(new_n510_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(KEYINPUT58), .C1(new_n762_), .C2(new_n758_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n559_), .A2(new_n783_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n758_), .A2(new_n762_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT58), .B1(new_n785_), .B2(new_n782_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n780_), .A2(new_n781_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n745_), .B1(new_n789_), .B2(new_n574_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n598_), .A2(new_n595_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(new_n334_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n738_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n787_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n573_), .B1(new_n796_), .B2(new_n781_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT59), .B(new_n793_), .C1(new_n797_), .C2(new_n745_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n423_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(G113gat), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT116), .B(new_n793_), .C1(new_n797_), .C2(new_n745_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n591_), .A2(new_n800_), .ZN(new_n805_));
  OAI22_X1  g604(.A1(new_n799_), .A2(new_n800_), .B1(new_n804_), .B2(new_n805_), .ZN(G1340gat));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT60), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n521_), .A2(KEYINPUT60), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n807_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n802_), .A2(new_n803_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n521_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n807_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT117), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n811_), .C1(new_n812_), .C2(new_n807_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1341gat));
  INV_X1    g616(.A(G127gat), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n802_), .A2(new_n803_), .A3(new_n818_), .A4(new_n573_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n574_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n818_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT118), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n823_), .B(new_n819_), .C1(new_n820_), .C2(new_n818_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1342gat));
  AOI21_X1  g624(.A(new_n623_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n826_));
  INV_X1    g625(.A(G134gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n589_), .A2(new_n827_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n826_), .A2(new_n827_), .B1(new_n804_), .B2(new_n828_), .ZN(G1343gat));
  NOR3_X1   g628(.A1(new_n790_), .A2(new_n331_), .A3(new_n792_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n591_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT119), .B(G141gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n578_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g634(.A1(new_n789_), .A2(new_n574_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n745_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n331_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n791_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT120), .B1(new_n840_), .B2(new_n574_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n830_), .A2(new_n842_), .A3(new_n573_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT61), .B(G155gat), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1346gat));
  INV_X1    g646(.A(G162gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n830_), .B2(new_n559_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n589_), .A2(new_n848_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n840_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT121), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1347gat));
  NOR2_X1   g655(.A1(new_n371_), .A2(new_n244_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n607_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n838_), .A2(new_n332_), .A3(new_n591_), .A4(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n283_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT122), .B1(new_n860_), .B2(G169gat), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(G169gat), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT62), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n867_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n865_), .B1(new_n869_), .B2(new_n870_), .ZN(G1348gat));
  NAND4_X1  g670(.A1(new_n838_), .A2(new_n332_), .A3(new_n578_), .A4(new_n859_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n282_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n790_), .A2(new_n281_), .ZN(new_n876_));
  INV_X1    g675(.A(G176gat), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n578_), .A4(new_n859_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n874_), .A2(new_n875_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n874_), .B2(new_n878_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1349gat));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n859_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n574_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n883_), .B(new_n298_), .C1(KEYINPUT124), .C2(G183gat), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(G183gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n883_), .B2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n882_), .B2(new_n623_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n589_), .A2(new_n299_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n882_), .B2(new_n889_), .ZN(G1351gat));
  NOR3_X1   g689(.A1(new_n790_), .A2(new_n331_), .A3(new_n858_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n591_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n578_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n896_));
  INV_X1    g695(.A(G211gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n573_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT125), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n891_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n897_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1354gat));
  NAND4_X1  g701(.A1(new_n838_), .A2(new_n839_), .A3(new_n589_), .A4(new_n857_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT127), .B(G218gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n623_), .A2(new_n906_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n905_), .A2(new_n906_), .B1(new_n891_), .B2(new_n907_), .ZN(G1355gat));
endmodule


