//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(KEYINPUT82), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n203_), .B1(new_n204_), .B2(KEYINPUT23), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT81), .B1(new_n207_), .B2(KEYINPUT26), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n206_), .B(new_n208_), .C1(new_n209_), .C2(KEYINPUT81), .ZN(new_n210_));
  NOR3_X1   g009(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n211_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n205_), .A2(new_n210_), .A3(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n202_), .A2(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n217_), .B(new_n219_), .C1(new_n204_), .C2(new_n218_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(G169gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n216_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G227gat), .A2(G233gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G15gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n224_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G71gat), .B(G99gat), .ZN(new_n228_));
  INV_X1    g027(.A(G43gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n227_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT84), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT85), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n237_), .B(KEYINPUT84), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n240_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n237_), .A2(KEYINPUT84), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(KEYINPUT84), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n241_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n242_), .B1(new_n248_), .B2(KEYINPUT85), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT31), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT86), .Z(new_n251_));
  NAND2_X1  g050(.A1(new_n236_), .A2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n250_), .A2(KEYINPUT86), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n234_), .A2(new_n253_), .A3(new_n235_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n257_), .B(KEYINPUT87), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G141gat), .B(G148gat), .Z(new_n267_));
  NAND3_X1  g066(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G141gat), .ZN(new_n271_));
  INV_X1    g070(.A(G148gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT89), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(KEYINPUT89), .ZN(new_n276_));
  OAI221_X1 g075(.A(new_n270_), .B1(KEYINPUT3), .B2(new_n273_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n259_), .A2(new_n262_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n266_), .A2(new_n267_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(KEYINPUT28), .ZN(new_n282_));
  XOR2_X1   g081(.A(G197gat), .B(G204gat), .Z(new_n283_));
  OR2_X1    g082(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n279_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT29), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n281_), .A2(KEYINPUT28), .ZN(new_n293_));
  OR3_X1    g092(.A1(new_n282_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n282_), .B2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(G78gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G106gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G22gat), .B(G50gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n294_), .A2(new_n295_), .A3(new_n301_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G8gat), .B(G36gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT18), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G64gat), .B(G92gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n214_), .A2(KEYINPUT93), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n214_), .A2(KEYINPUT93), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT94), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n313_), .A2(KEYINPUT94), .A3(new_n314_), .A4(new_n315_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n318_), .A2(new_n319_), .B1(new_n205_), .B2(new_n217_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n219_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n202_), .B(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n323_), .B2(KEYINPUT23), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n215_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n206_), .A2(KEYINPUT91), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n206_), .A2(KEYINPUT91), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n209_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT92), .B1(new_n332_), .B2(new_n325_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n320_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n290_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n224_), .B2(new_n289_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n335_), .A2(new_n336_), .A3(new_n339_), .A4(new_n341_), .ZN(new_n342_));
  AOI211_X1 g141(.A(new_n289_), .B(new_n320_), .C1(new_n331_), .C2(new_n333_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n339_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT95), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n320_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n327_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n332_), .A2(new_n325_), .A3(KEYINPUT92), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n224_), .B2(new_n289_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n350_), .A2(new_n289_), .B1(new_n351_), .B2(KEYINPUT90), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(KEYINPUT90), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n339_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n310_), .B1(new_n346_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(KEYINPUT90), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n290_), .B2(new_n334_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n338_), .B1(new_n358_), .B2(new_n353_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(new_n309_), .A3(new_n342_), .A4(new_n345_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n291_), .A2(new_n249_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n279_), .A2(new_n248_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n291_), .A2(new_n249_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT97), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n291_), .A2(new_n249_), .A3(KEYINPUT97), .A4(new_n372_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n248_), .A2(KEYINPUT85), .ZN(new_n379_));
  INV_X1    g178(.A(new_n242_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n364_), .B(KEYINPUT4), .C1(new_n381_), .C2(new_n279_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n362_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n371_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n356_), .A2(new_n360_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n363_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT98), .B1(new_n378_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n370_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n382_), .A2(new_n363_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT98), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n377_), .A3(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .A4(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n385_), .B1(new_n386_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n390_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n392_), .B1(new_n391_), .B2(new_n377_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT100), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(KEYINPUT33), .A4(new_n389_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT100), .B1(new_n394_), .B2(new_n386_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n370_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n394_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n359_), .A2(KEYINPUT101), .A3(new_n342_), .A4(new_n345_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n326_), .A2(new_n330_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n347_), .A2(new_n290_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n339_), .B1(new_n407_), .B2(new_n341_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT102), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n309_), .A2(KEYINPUT32), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n352_), .A2(new_n339_), .A3(new_n354_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n405_), .A2(new_n409_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n346_), .A2(new_n355_), .A3(KEYINPUT101), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n404_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n305_), .B1(new_n402_), .B2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n409_), .A2(new_n412_), .ZN(new_n418_));
  OAI211_X1 g217(.A(KEYINPUT27), .B(new_n360_), .C1(new_n418_), .C2(new_n309_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT27), .B1(new_n356_), .B2(new_n360_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(KEYINPUT103), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT103), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n422_), .B(KEYINPUT27), .C1(new_n356_), .C2(new_n360_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n403_), .A2(new_n394_), .A3(new_n305_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n255_), .B1(new_n417_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n424_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n255_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n404_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n305_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G29gat), .B(G36gat), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n434_), .A2(KEYINPUT75), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(KEYINPUT75), .ZN(new_n436_));
  XOR2_X1   g235(.A(G43gat), .B(G50gat), .Z(new_n437_));
  OR3_X1    g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT15), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G22gat), .ZN(new_n442_));
  INV_X1    g241(.A(G1gat), .ZN(new_n443_));
  INV_X1    g242(.A(G8gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT14), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G8gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n441_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n440_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n440_), .B(new_n451_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(G229gat), .A3(G233gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G113gat), .B(G141gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G169gat), .B(G197gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT80), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(KEYINPUT80), .A3(new_n462_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G231gat), .A2(G233gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n448_), .B(new_n468_), .Z(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G64gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G71gat), .B(G78gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT11), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n473_));
  INV_X1    g272(.A(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n469_), .B(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n478_), .A2(KEYINPUT68), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(KEYINPUT68), .ZN(new_n480_));
  XOR2_X1   g279(.A(G127gat), .B(G155gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G183gat), .B(G211gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(KEYINPUT17), .Z(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n480_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT78), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n478_), .A2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT79), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(KEYINPUT79), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT9), .ZN(new_n495_));
  AND2_X1   g294(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT65), .B(G92gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  AND2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(KEYINPUT9), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT6), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(G99gat), .A3(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n504_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519_));
  INV_X1    g318(.A(G99gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n506_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n511_), .B1(G99gat), .B2(G106gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n509_), .A2(KEYINPUT6), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n518_), .B(new_n521_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT66), .B1(new_n502_), .B2(new_n501_), .ZN(new_n525_));
  INV_X1    g324(.A(G85gat), .ZN(new_n526_));
  INV_X1    g325(.A(G92gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AND4_X1   g330(.A1(new_n517_), .A2(new_n524_), .A3(new_n525_), .A4(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n525_), .A2(new_n531_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n517_), .B1(new_n533_), .B2(new_n524_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n516_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n441_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(KEYINPUT67), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n510_), .A2(new_n512_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n521_), .A2(new_n518_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n525_), .A2(new_n531_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT8), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n533_), .A2(new_n517_), .A3(new_n524_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n516_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n537_), .A2(new_n440_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n536_), .B(new_n547_), .C1(KEYINPUT35), .C2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT36), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n555_), .A2(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n552_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT37), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n558_), .A2(new_n563_), .A3(new_n560_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n494_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n477_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n544_), .B2(new_n516_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n477_), .A2(KEYINPUT68), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT68), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n572_), .B(new_n472_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n537_), .A2(new_n546_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n537_), .B2(new_n546_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT12), .ZN(new_n580_));
  INV_X1    g379(.A(new_n574_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n514_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n582_));
  AOI211_X1 g381(.A(KEYINPUT67), .B(new_n582_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n545_), .B1(new_n544_), .B2(new_n516_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT70), .B1(new_n585_), .B2(new_n567_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n570_), .B(new_n577_), .C1(new_n580_), .C2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT69), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n575_), .B(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n576_), .B1(new_n590_), .B2(new_n585_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G176gat), .B(G204gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT72), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT73), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n593_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n588_), .A2(new_n591_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(KEYINPUT13), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(KEYINPUT13), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n601_), .B(new_n602_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n601_), .A2(new_n602_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n606_), .B1(new_n607_), .B2(new_n605_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n566_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n433_), .A2(new_n467_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT104), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n443_), .A3(new_n404_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n561_), .B(KEYINPUT105), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n467_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n494_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT106), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n443_), .B1(new_n622_), .B2(new_n404_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n615_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n614_), .B2(new_n613_), .ZN(G1324gat));
  OAI21_X1  g424(.A(G8gat), .B1(new_n621_), .B2(new_n428_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT39), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n428_), .A2(G8gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT107), .B1(new_n612_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n611_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT104), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n611_), .A2(new_n632_), .ZN(new_n633_));
  AND4_X1   g432(.A1(KEYINPUT107), .A2(new_n631_), .A3(new_n633_), .A4(new_n628_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n627_), .B1(new_n629_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n627_), .B(KEYINPUT40), .C1(new_n629_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  OR3_X1    g438(.A1(new_n611_), .A2(G15gat), .A3(new_n255_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n622_), .A2(new_n429_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n641_), .B2(G15gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  INV_X1    g443(.A(G22gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n630_), .A2(new_n645_), .A3(new_n305_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n622_), .A2(new_n305_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(G22gat), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT42), .B(new_n645_), .C1(new_n622_), .C2(new_n305_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1327gat));
  INV_X1    g450(.A(new_n494_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n561_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n433_), .A2(new_n467_), .A3(new_n608_), .A4(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G29gat), .B1(new_n655_), .B2(new_n404_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n619_), .A2(new_n652_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n562_), .A2(new_n564_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n433_), .B2(new_n660_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT43), .B(new_n659_), .C1(new_n427_), .C2(new_n432_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT44), .B(new_n657_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n404_), .A2(G29gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n656_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n424_), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n654_), .A2(G36gat), .A3(new_n428_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(KEYINPUT46), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  NAND4_X1  g478(.A1(new_n665_), .A2(G43gat), .A3(new_n429_), .A4(new_n666_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n229_), .B1(new_n654_), .B2(new_n255_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g482(.A1(new_n654_), .A2(G50gat), .A3(new_n431_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n665_), .A2(new_n305_), .A3(new_n666_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(G50gat), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT108), .B(new_n684_), .C1(new_n685_), .C2(G50gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1331gat));
  NOR3_X1   g489(.A1(new_n608_), .A2(new_n467_), .A3(new_n494_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n618_), .A2(G57gat), .A3(new_n404_), .A4(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT111), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n467_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n609_), .A3(new_n565_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n430_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n699_), .B1(new_n698_), .B2(new_n697_), .ZN(new_n700_));
  INV_X1    g499(.A(G57gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n693_), .B1(new_n700_), .B2(new_n701_), .ZN(G1332gat));
  NAND3_X1  g501(.A1(new_n618_), .A2(new_n424_), .A3(new_n691_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G64gat), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT48), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT48), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n428_), .A2(G64gat), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n705_), .A2(new_n706_), .B1(new_n697_), .B2(new_n707_), .ZN(G1333gat));
  OR3_X1    g507(.A1(new_n697_), .A2(G71gat), .A3(new_n255_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n618_), .A2(new_n429_), .A3(new_n691_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(G71gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n711_), .B2(G71gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n714_), .A2(new_n710_), .A3(new_n715_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n709_), .A2(new_n716_), .A3(new_n717_), .ZN(G1334gat));
  NAND3_X1  g517(.A1(new_n618_), .A2(new_n305_), .A3(new_n691_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G78gat), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT50), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT50), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n431_), .A2(G78gat), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n721_), .A2(new_n722_), .B1(new_n697_), .B2(new_n723_), .ZN(G1335gat));
  OR2_X1    g523(.A1(new_n661_), .A2(new_n662_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n608_), .A2(new_n467_), .A3(new_n652_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n430_), .A2(new_n498_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n608_), .A2(new_n652_), .A3(new_n561_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n696_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n526_), .B1(new_n732_), .B2(new_n430_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT113), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n730_), .A2(new_n736_), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1336gat));
  NOR2_X1   g537(.A1(new_n428_), .A2(new_n499_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n728_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n527_), .B1(new_n732_), .B2(new_n428_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT114), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1337gat));
  OAI21_X1  g545(.A(G99gat), .B1(new_n727_), .B2(new_n255_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n429_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n732_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n747_), .B(new_n751_), .C1(new_n732_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  OAI211_X1 g552(.A(new_n726_), .B(new_n305_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G106gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n305_), .A2(new_n506_), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n756_), .A2(new_n757_), .B1(new_n732_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g559(.A(new_n467_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n565_), .A2(new_n608_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT115), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n565_), .A2(new_n608_), .A3(new_n764_), .A4(new_n761_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(KEYINPUT54), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(KEYINPUT115), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n561_), .A2(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n449_), .A2(new_n452_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT118), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT118), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n450_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n459_), .B1(new_n454_), .B2(new_n450_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n462_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n607_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n467_), .A2(new_n601_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n587_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n579_), .B1(new_n578_), .B2(KEYINPUT12), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n585_), .A2(KEYINPUT70), .A3(new_n567_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n569_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n577_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n590_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n784_), .A2(new_n785_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n590_), .A3(new_n570_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n576_), .B1(new_n792_), .B2(KEYINPUT116), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n788_), .B1(new_n790_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n781_), .B1(new_n794_), .B2(new_n598_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n796_));
  INV_X1    g595(.A(new_n576_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n790_), .ZN(new_n798_));
  AND4_X1   g597(.A1(KEYINPUT55), .A2(new_n791_), .A3(new_n570_), .A4(new_n577_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT55), .B1(new_n786_), .B2(new_n577_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n599_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n780_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n779_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n780_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n599_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n781_), .B(new_n598_), .C1(new_n798_), .C2(new_n801_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(KEYINPUT117), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n770_), .B1(new_n806_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n777_), .A2(new_n600_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT120), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n659_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n795_), .A2(new_n803_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT58), .A4(new_n813_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n561_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n778_), .B1(new_n810_), .B2(KEYINPUT117), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n812_), .B(new_n821_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n769_), .B1(new_n827_), .B2(new_n494_), .ZN(new_n828_));
  NOR4_X1   g627(.A1(new_n424_), .A2(new_n255_), .A3(new_n430_), .A4(new_n305_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n467_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(KEYINPUT59), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n761_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n833_), .B1(new_n837_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(KEYINPUT60), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(KEYINPUT121), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n831_), .B(new_n842_), .C1(KEYINPUT121), .C2(new_n840_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n608_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n839_), .ZN(G1341gat));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n831_), .A2(new_n846_), .A3(new_n652_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n494_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n846_), .ZN(G1342gat));
  NOR3_X1   g648(.A1(new_n828_), .A2(new_n616_), .A3(new_n830_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT122), .B1(new_n850_), .B2(G134gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n834_), .A2(new_n836_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n659_), .A2(new_n853_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n854_), .A2(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n812_), .A2(new_n821_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n810_), .A2(KEYINPUT117), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n824_), .A3(new_n779_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n826_), .B1(new_n861_), .B2(new_n561_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n494_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n769_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n429_), .A2(new_n431_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n404_), .A3(new_n428_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT123), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n828_), .A2(new_n870_), .A3(new_n867_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n467_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G141gat), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n271_), .B(new_n467_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1344gat));
  OAI21_X1  g674(.A(new_n609_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G148gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n272_), .B(new_n609_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1345gat));
  OAI21_X1  g678(.A(new_n652_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n881_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n652_), .B(new_n883_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n617_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n865_), .A2(KEYINPUT123), .A3(new_n868_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n870_), .B1(new_n828_), .B2(new_n867_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n659_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n886_), .B2(new_n890_), .ZN(G1347gat));
  NAND3_X1  g690(.A1(new_n424_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT124), .ZN(new_n893_));
  NOR4_X1   g692(.A1(new_n828_), .A2(new_n305_), .A3(new_n761_), .A4(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(G169gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(new_n897_), .A3(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n898_), .B(new_n899_), .C1(new_n894_), .C2(new_n896_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n894_), .A2(new_n311_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(G1348gat));
  NOR3_X1   g703(.A1(new_n828_), .A2(new_n305_), .A3(new_n893_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n609_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g706(.A(G183gat), .B1(new_n905_), .B2(new_n652_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n328_), .A2(new_n329_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n905_), .A2(new_n652_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1350gat));
  NAND3_X1  g710(.A1(new_n905_), .A2(new_n209_), .A3(new_n617_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n905_), .A2(new_n660_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n207_), .ZN(G1351gat));
  NOR4_X1   g713(.A1(new_n428_), .A2(new_n429_), .A3(new_n404_), .A4(new_n431_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n865_), .A2(G197gat), .A3(new_n467_), .A4(new_n915_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n916_), .A2(KEYINPUT126), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(KEYINPUT126), .ZN(new_n918_));
  INV_X1    g717(.A(G197gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n865_), .A2(new_n915_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n761_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n917_), .A2(new_n918_), .A3(new_n921_), .ZN(G1352gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n608_), .ZN(new_n923_));
  INV_X1    g722(.A(G204gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1353gat));
  OR2_X1    g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n920_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n652_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n920_), .A2(new_n494_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT63), .B(G211gat), .Z(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(G1354gat));
  AOI21_X1  g730(.A(G218gat), .B1(new_n927_), .B2(new_n617_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n660_), .A2(G218gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT127), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n927_), .B2(new_n934_), .ZN(G1355gat));
endmodule


