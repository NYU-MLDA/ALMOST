//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT95), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  OR3_X1    g004(.A1(new_n205_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT93), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(G204gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n203_), .A2(KEYINPUT95), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT91), .ZN(new_n215_));
  OR3_X1    g014(.A1(new_n205_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT21), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT92), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n206_), .A2(new_n209_), .A3(new_n219_), .A4(new_n210_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT92), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n215_), .A2(new_n216_), .A3(new_n221_), .A4(KEYINPUT21), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n218_), .A2(new_n220_), .A3(new_n202_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT94), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n220_), .A2(new_n202_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT94), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n222_), .A4(new_n218_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n214_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT24), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT23), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G183gat), .A3(G190gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n234_), .A2(KEYINPUT24), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n237_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(KEYINPUT83), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n238_), .B2(KEYINPUT23), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(G183gat), .B2(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n235_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G169gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n233_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n244_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n228_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT19), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n235_), .B1(new_n242_), .B2(new_n259_), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n232_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT22), .B1(new_n232_), .B2(KEYINPUT85), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n261_), .A2(new_n233_), .A3(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n243_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n248_), .A2(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(KEYINPUT84), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n237_), .B1(new_n266_), .B2(KEYINPUT84), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT99), .B1(new_n258_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n224_), .A2(new_n227_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n213_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n256_), .B1(new_n228_), .B2(new_n253_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT99), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .A4(KEYINPUT20), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n228_), .A2(new_n269_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n253_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n256_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n271_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT18), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n271_), .A2(new_n282_), .A3(new_n278_), .A4(new_n287_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n254_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n256_), .B1(new_n294_), .B2(new_n270_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n228_), .A2(new_n253_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(KEYINPUT20), .A3(new_n257_), .A4(new_n279_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n288_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT27), .A3(new_n290_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT102), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n299_), .A2(new_n290_), .A3(KEYINPUT102), .A4(KEYINPUT27), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n293_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n269_), .A2(KEYINPUT30), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n269_), .A2(KEYINPUT30), .ZN(new_n308_));
  OAI21_X1  g107(.A(G99gat), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  INV_X1    g109(.A(G99gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(new_n306_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n305_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G227gat), .A2(G233gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(G15gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G71gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT86), .B(G43gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT87), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n318_), .B(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322_));
  XOR2_X1   g121(.A(G113gat), .B(G120gat), .Z(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n321_), .B(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n314_), .A2(new_n315_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n315_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(new_n313_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT89), .ZN(new_n339_));
  INV_X1    g138(.A(G141gat), .ZN(new_n340_));
  INV_X1    g139(.A(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT88), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n343_), .A2(new_n340_), .A3(new_n341_), .A4(KEYINPUT88), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n345_), .B(new_n346_), .C1(new_n337_), .C2(new_n336_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n334_), .B(new_n335_), .C1(new_n339_), .C2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n333_), .B1(KEYINPUT1), .B2(new_n335_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(KEYINPUT1), .B2(new_n335_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n336_), .A3(new_n342_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(KEYINPUT100), .A3(new_n324_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n351_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT100), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n325_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n332_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n325_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G85gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n357_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n369_), .B1(new_n372_), .B2(new_n364_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT101), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(KEYINPUT101), .B(new_n369_), .C1(new_n372_), .C2(new_n364_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n331_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT98), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT90), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n352_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n228_), .B2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n381_), .B1(new_n354_), .B2(KEYINPUT29), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n273_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT28), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n352_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT28), .B1(new_n354_), .B2(KEYINPUT29), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G22gat), .B(G50gat), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n388_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n389_), .B(new_n397_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n398_), .A2(new_n399_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n379_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n398_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT97), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n397_), .A2(new_n389_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n398_), .A2(new_n399_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT98), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n397_), .B1(new_n403_), .B2(new_n389_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n304_), .A2(new_n378_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n359_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(new_n370_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT33), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n371_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n363_), .A2(KEYINPUT33), .A3(new_n365_), .A4(new_n370_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n289_), .A3(new_n290_), .A4(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n298_), .A2(KEYINPUT32), .A3(new_n287_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n287_), .A2(KEYINPUT32), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n422_), .B2(new_n283_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n377_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n409_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n411_), .A2(new_n377_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n304_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n331_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n412_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G229gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G1gat), .B(G8gat), .Z(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G15gat), .B(G22gat), .Z(new_n435_));
  NAND2_X1  g234(.A1(G1gat), .A2(G8gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT14), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT78), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT79), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n437_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n440_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n434_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n443_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n442_), .B1(new_n441_), .B2(new_n437_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT79), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n433_), .A3(new_n444_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G29gat), .B(G36gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G43gat), .B(G50gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n447_), .A2(new_n451_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n432_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n455_), .B(KEYINPUT15), .ZN(new_n459_));
  INV_X1    g258(.A(new_n451_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n433_), .B1(new_n450_), .B2(new_n444_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n447_), .A2(new_n451_), .A3(new_n455_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n431_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n458_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G113gat), .B(G141gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G169gat), .B(G197gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n466_), .B(new_n467_), .Z(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n458_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT82), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(KEYINPUT82), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n430_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT9), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n477_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT65), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n478_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n478_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n481_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(KEYINPUT65), .A3(new_n484_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT64), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT6), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n502_), .A2(new_n504_), .A3(KEYINPUT66), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT66), .B1(new_n502_), .B2(new_n504_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n500_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n491_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(new_n504_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT67), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT68), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(new_n311_), .A3(new_n495_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT68), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n512_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n502_), .A2(new_n504_), .A3(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n511_), .A2(new_n515_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n479_), .A2(new_n480_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n509_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n509_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n505_), .A2(new_n506_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n513_), .A2(new_n514_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n508_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G71gat), .B(G78gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(KEYINPUT11), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(KEYINPUT11), .ZN(new_n533_));
  INV_X1    g332(.A(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n530_), .A2(KEYINPUT11), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n529_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n537_), .B(new_n508_), .C1(new_n524_), .C2(new_n528_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G230gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n542_), .B(new_n544_), .C1(new_n540_), .C2(new_n539_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT12), .B1(new_n529_), .B2(new_n538_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n538_), .A2(KEYINPUT12), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT70), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n494_), .A2(new_n499_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n526_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n550_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n491_), .A2(new_n507_), .A3(KEYINPUT70), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n524_), .A2(new_n528_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n549_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n547_), .A2(new_n560_), .A3(new_n543_), .A4(new_n541_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n545_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n545_), .A2(new_n561_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(KEYINPUT13), .A3(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT80), .Z(new_n577_));
  NOR3_X1   g376(.A1(new_n460_), .A2(new_n461_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n582_), .A3(new_n538_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n537_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n583_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT81), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n594_));
  INV_X1    g393(.A(new_n583_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n590_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G190gat), .B(G218gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT73), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT75), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n522_), .A2(new_n523_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT8), .ZN(new_n613_));
  INV_X1    g412(.A(new_n528_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n613_), .A2(new_n614_), .B1(new_n491_), .B2(new_n507_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n611_), .B1(new_n615_), .B2(new_n455_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n608_), .A2(new_n609_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n556_), .B(new_n557_), .C1(new_n524_), .C2(new_n528_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n459_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n616_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n605_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n616_), .A2(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n617_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n616_), .A2(new_n620_), .A3(new_n618_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n603_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n623_), .A2(new_n629_), .A3(KEYINPUT37), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT77), .B1(new_n621_), .B2(new_n622_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n625_), .A2(new_n632_), .A3(new_n626_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n633_), .A3(new_n605_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(new_n629_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n635_), .B2(KEYINPUT37), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n475_), .A2(new_n575_), .A3(new_n599_), .A4(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G1gat), .A3(new_n377_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n430_), .A2(new_n635_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n472_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n574_), .A2(new_n643_), .A3(new_n598_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n377_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n639_), .A2(new_n640_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n641_), .A2(new_n647_), .A3(new_n648_), .ZN(G1324gat));
  AND3_X1   g448(.A1(new_n293_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n638_), .A2(G8gat), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n645_), .A2(new_n304_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G8gat), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n653_), .A2(KEYINPUT39), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(KEYINPUT39), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n646_), .B2(new_n429_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n638_), .A2(G15gat), .A3(new_n429_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1326gat));
  OR3_X1    g461(.A1(new_n638_), .A2(G22gat), .A3(new_n425_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n645_), .A2(new_n411_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G22gat), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(KEYINPUT42), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(KEYINPUT42), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(G1327gat));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n430_), .B2(new_n637_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  AOI22_X1  g471(.A1(new_n408_), .A2(new_n410_), .B1(new_n376_), .B2(new_n375_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n650_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n331_), .B1(new_n674_), .B2(new_n426_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n672_), .B(new_n636_), .C1(new_n675_), .C2(new_n412_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n574_), .A2(new_n643_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n598_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT44), .B1(new_n677_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n682_), .B(new_n679_), .C1(new_n671_), .C2(new_n676_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n681_), .A2(new_n683_), .A3(new_n377_), .ZN(new_n684_));
  INV_X1    g483(.A(G29gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n635_), .A2(new_n598_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n574_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n475_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n377_), .A2(G29gat), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT105), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n684_), .A2(new_n685_), .B1(new_n688_), .B2(new_n690_), .ZN(G1328gat));
  NOR3_X1   g490(.A1(new_n688_), .A2(G36gat), .A3(new_n650_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n677_), .A2(new_n680_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n682_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n677_), .A2(KEYINPUT44), .A3(new_n680_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n304_), .A4(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n681_), .A2(new_n683_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n701_), .B2(new_n304_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n694_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT46), .B(new_n694_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  NAND3_X1  g506(.A1(new_n701_), .A2(G43gat), .A3(new_n331_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n688_), .A2(new_n429_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(G43gat), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(G1330gat));
  OR3_X1    g511(.A1(new_n688_), .A2(G50gat), .A3(new_n425_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n701_), .A2(new_n714_), .A3(new_n411_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G50gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n701_), .B2(new_n411_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1331gat));
  NAND4_X1  g517(.A1(new_n474_), .A2(new_n473_), .A3(new_n593_), .A4(new_n597_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n575_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n642_), .A2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n377_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n430_), .A2(new_n472_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(new_n574_), .A3(new_n599_), .A4(new_n637_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n377_), .A2(G57gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(G1332gat));
  OAI21_X1  g525(.A(G64gat), .B1(new_n721_), .B2(new_n650_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT48), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n650_), .A2(G64gat), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT109), .Z(new_n730_));
  OAI21_X1  g529(.A(new_n728_), .B1(new_n724_), .B2(new_n730_), .ZN(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n721_), .B2(new_n429_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT49), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n429_), .A2(G71gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n724_), .B2(new_n734_), .ZN(G1334gat));
  OAI21_X1  g534(.A(G78gat), .B1(new_n721_), .B2(new_n425_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT50), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n425_), .A2(G78gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n724_), .B2(new_n738_), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n575_), .A2(new_n686_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n723_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n476_), .B1(new_n741_), .B2(new_n377_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT110), .Z(new_n743_));
  NOR3_X1   g542(.A1(new_n575_), .A2(new_n472_), .A3(new_n599_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n677_), .A2(new_n744_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n745_), .A2(new_n476_), .A3(new_n377_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n745_), .B2(new_n650_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n304_), .A2(new_n477_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n741_), .B2(new_n749_), .ZN(G1337gat));
  OAI21_X1  g549(.A(G99gat), .B1(new_n745_), .B2(new_n429_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n331_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n741_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g553(.A1(new_n741_), .A2(new_n425_), .A3(new_n499_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n756_));
  INV_X1    g555(.A(new_n745_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n411_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n758_), .B2(G106gat), .ZN(new_n759_));
  INV_X1    g558(.A(new_n756_), .ZN(new_n760_));
  AOI211_X1 g559(.A(new_n495_), .B(new_n760_), .C1(new_n757_), .C2(new_n411_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n755_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n755_), .C1(new_n759_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  INV_X1    g565(.A(KEYINPUT59), .ZN(new_n767_));
  NOR4_X1   g566(.A1(new_n304_), .A2(new_n411_), .A3(new_n429_), .A4(new_n377_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n472_), .A2(new_n569_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n541_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n619_), .B2(new_n549_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n543_), .B1(new_n772_), .B2(new_n547_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n561_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n560_), .A2(new_n541_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n544_), .B1(new_n776_), .B2(new_n546_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n491_), .A2(new_n507_), .A3(KEYINPUT70), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT70), .B1(new_n491_), .B2(new_n507_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n613_), .A2(new_n614_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n548_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NOR4_X1   g581(.A1(new_n782_), .A2(new_n546_), .A3(new_n544_), .A4(new_n771_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n777_), .A2(new_n783_), .A3(KEYINPUT55), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n775_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n566_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n787_), .B(new_n568_), .C1(new_n775_), .C2(new_n784_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n770_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n431_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n462_), .A2(new_n463_), .A3(new_n432_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n469_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n471_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n569_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n568_), .B1(new_n545_), .B2(new_n561_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n790_), .B(new_n794_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n790_), .B1(new_n570_), .B2(new_n794_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n789_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n635_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT57), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n635_), .C1(new_n789_), .C2(new_n800_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n794_), .A2(new_n569_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n783_), .B1(KEYINPUT55), .B2(new_n777_), .ZN(new_n808_));
  NOR4_X1   g607(.A1(new_n776_), .A2(new_n774_), .A3(new_n544_), .A4(new_n546_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n566_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n787_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n807_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n636_), .B1(new_n813_), .B2(KEYINPUT58), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(KEYINPUT58), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT114), .B(new_n636_), .C1(new_n813_), .C2(KEYINPUT58), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n599_), .B1(new_n806_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  OR3_X1    g620(.A1(new_n719_), .A2(new_n574_), .A3(KEYINPUT112), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT112), .B1(new_n719_), .B2(new_n574_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n821_), .B1(new_n824_), .B2(new_n637_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT54), .B(new_n636_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n767_), .B(new_n768_), .C1(new_n820_), .C2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n768_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n818_), .A2(new_n817_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n807_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT114), .B1(new_n834_), .B2(new_n636_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n830_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n769_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT113), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n797_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n802_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n804_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n801_), .A2(KEYINPUT57), .A3(new_n802_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT115), .B1(new_n836_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n806_), .A2(new_n819_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n598_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n827_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n829_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n828_), .B1(new_n850_), .B2(new_n767_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n474_), .A2(new_n473_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n828_), .B(KEYINPUT116), .C1(new_n850_), .C2(new_n767_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G113gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n850_), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n858_), .A2(G113gat), .A3(new_n643_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1340gat));
  INV_X1    g659(.A(G120gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n850_), .B(new_n862_), .C1(KEYINPUT60), .C2(new_n861_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n851_), .A2(new_n575_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n865_), .B2(new_n861_), .ZN(G1341gat));
  AND2_X1   g665(.A1(new_n853_), .A2(new_n855_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT118), .B(G127gat), .Z(new_n868_));
  NOR2_X1   g667(.A1(new_n598_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n858_), .B2(new_n598_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT117), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n873_), .B(new_n870_), .C1(new_n858_), .C2(new_n598_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n867_), .A2(new_n869_), .B1(new_n872_), .B2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n850_), .B2(new_n635_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT119), .B(G134gat), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n637_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n867_), .B2(new_n878_), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n848_), .A2(new_n849_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n304_), .A2(new_n425_), .A3(new_n377_), .A4(new_n331_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(KEYINPUT120), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(KEYINPUT120), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n472_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G141gat), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n340_), .B(new_n472_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1344gat));
  OAI21_X1  g687(.A(new_n574_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G148gat), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n341_), .B(new_n574_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1345gat));
  OAI21_X1  g691(.A(new_n599_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n894_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n599_), .B(new_n896_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1346gat));
  INV_X1    g697(.A(new_n884_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n882_), .A2(KEYINPUT120), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n637_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(G162gat), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n883_), .A2(new_n884_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n635_), .A2(new_n902_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n901_), .A2(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(G1347gat));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n820_), .A2(new_n827_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n650_), .A2(new_n378_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT121), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n411_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n643_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n906_), .B1(new_n912_), .B2(new_n232_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n251_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT62), .B(G169gat), .C1(new_n911_), .C2(new_n643_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  OAI21_X1  g715(.A(new_n233_), .B1(new_n911_), .B2(new_n575_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n918_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n411_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n909_), .A2(new_n233_), .A3(new_n575_), .ZN(new_n922_));
  AOI22_X1  g721(.A1(new_n919_), .A2(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1349gat));
  NOR3_X1   g722(.A1(new_n911_), .A2(new_n229_), .A3(new_n598_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT123), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n909_), .A2(new_n598_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G183gat), .B1(new_n921_), .B2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n911_), .B2(new_n637_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n635_), .A2(new_n230_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n911_), .B2(new_n930_), .ZN(G1351gat));
  NAND2_X1  g730(.A1(new_n673_), .A2(new_n429_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n304_), .B1(new_n932_), .B2(KEYINPUT124), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n933_), .B1(KEYINPUT124), .B2(new_n932_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n880_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n472_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n205_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(KEYINPUT126), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(new_n939_), .A3(new_n205_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n936_), .B2(new_n205_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n935_), .A2(new_n942_), .A3(G197gat), .A4(new_n472_), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n938_), .A2(new_n940_), .B1(new_n941_), .B2(new_n943_), .ZN(G1352gat));
  NAND2_X1  g743(.A1(new_n935_), .A2(new_n574_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g745(.A1(new_n935_), .A2(new_n599_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  AND2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n950_), .B1(new_n947_), .B2(new_n948_), .ZN(G1354gat));
  NAND2_X1  g750(.A1(new_n935_), .A2(new_n635_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT127), .B(G218gat), .Z(new_n953_));
  NOR2_X1   g752(.A1(new_n637_), .A2(new_n953_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n952_), .A2(new_n953_), .B1(new_n935_), .B2(new_n954_), .ZN(G1355gat));
endmodule


