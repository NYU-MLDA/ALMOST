//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n208_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G85gat), .B(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  OR2_X1    g020(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n224_), .B2(KEYINPUT9), .ZN(new_n225_));
  AND2_X1   g024(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(G85gat), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT9), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT66), .A3(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n225_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT10), .B(G99gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n207_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n217_), .A2(new_n219_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G29gat), .B(G36gat), .Z(new_n244_));
  XOR2_X1   g043(.A(G43gat), .B(G50gat), .Z(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT15), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n244_), .B(new_n245_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT15), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n212_), .A2(new_n208_), .ZN(new_n252_));
  AOI211_X1 g051(.A(KEYINPUT8), .B(new_n214_), .C1(new_n252_), .C2(new_n207_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n218_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n228_), .A2(new_n229_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n233_), .B1(new_n256_), .B2(new_n220_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n239_), .B1(new_n257_), .B2(new_n230_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n243_), .A2(new_n251_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n241_), .A2(new_n248_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT73), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G232gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT35), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n260_), .A2(KEYINPUT73), .A3(new_n261_), .A4(new_n265_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G190gat), .B(G218gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(G134gat), .B(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT36), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n202_), .B1(new_n278_), .B2(KEYINPUT75), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT36), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT74), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n272_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT75), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n283_), .B(new_n284_), .C1(new_n272_), .C2(new_n277_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n279_), .A2(new_n285_), .A3(KEYINPUT76), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT76), .B1(new_n279_), .B2(new_n285_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n277_), .B1(new_n272_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n288_), .B2(new_n272_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n283_), .ZN(new_n291_));
  OAI22_X1  g090(.A1(new_n286_), .A2(new_n287_), .B1(KEYINPUT37), .B2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT78), .B(G1gat), .Z(new_n293_));
  INV_X1    g092(.A(G8gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT79), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n302_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G71gat), .B(G78gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G57gat), .B(G64gat), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(KEYINPUT11), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(KEYINPUT11), .B2(new_n307_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n306_), .A3(KEYINPUT11), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n305_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G127gat), .B(G155gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G183gat), .B(G211gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT17), .Z(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(KEYINPUT81), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(KEYINPUT17), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n319_), .B1(new_n312_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT81), .B1(new_n312_), .B2(new_n318_), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n292_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT83), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT13), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n311_), .A2(KEYINPUT12), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n243_), .A2(new_n333_), .A3(new_n259_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n309_), .A2(new_n310_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n241_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n217_), .A2(new_n219_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n235_), .A2(new_n240_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT12), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n311_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT12), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT68), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n334_), .B(new_n338_), .C1(new_n343_), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT69), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n241_), .A2(new_n337_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n336_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n342_), .B1(new_n341_), .B2(KEYINPUT12), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n344_), .A2(KEYINPUT68), .A3(new_n345_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT69), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n334_), .A4(new_n338_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n348_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G120gat), .B(G148gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(G176gat), .B(G204gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n348_), .A2(new_n351_), .A3(new_n356_), .A4(new_n362_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n365_), .A2(KEYINPUT71), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(KEYINPUT71), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n331_), .B(new_n364_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n365_), .B(KEYINPUT71), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n331_), .B1(new_n370_), .B2(new_n364_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n330_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT72), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(KEYINPUT13), .A3(new_n368_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(G176gat), .B1(KEYINPUT90), .B2(KEYINPUT22), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G169gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT23), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(G183gat), .A3(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n378_), .A2(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G183gat), .ZN(new_n395_));
  INV_X1    g194(.A(G183gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT25), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n393_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n393_), .B1(new_n396_), .B2(KEYINPUT25), .ZN(new_n399_));
  INV_X1    g198(.A(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT26), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT26), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G190gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n392_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n382_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n380_), .A2(KEYINPUT89), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n379_), .A2(new_n408_), .A3(KEYINPUT23), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n387_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT91), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n411_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(G15gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT30), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n419_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(KEYINPUT92), .A3(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G127gat), .B(G134gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n423_), .A2(new_n424_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT31), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n427_), .A2(KEYINPUT31), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT92), .B1(new_n420_), .B2(new_n421_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n430_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n437_));
  INV_X1    g236(.A(G141gat), .ZN(new_n438_));
  INV_X1    g237(.A(G148gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n438_), .A2(new_n439_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n441_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT1), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n447_), .A2(new_n454_), .A3(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n456_), .A3(KEYINPUT100), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n423_), .B(new_n424_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n446_), .A2(new_n449_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n427_), .A3(KEYINPUT100), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n436_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n460_), .A2(new_n458_), .A3(KEYINPUT4), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n435_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n459_), .A2(new_n461_), .A3(new_n434_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT101), .B(G85gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT0), .B(G57gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n464_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n433_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n450_), .A2(new_n456_), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n475_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT28), .B1(new_n475_), .B2(KEYINPUT29), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G22gat), .B(G50gat), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484_));
  OAI21_X1  g283(.A(G228gat), .B1(new_n484_), .B2(G233gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n484_), .B2(G233gat), .ZN(new_n486_));
  INV_X1    g285(.A(G211gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(G218gat), .ZN(new_n488_));
  INV_X1    g287(.A(G218gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(G211gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT96), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT95), .ZN(new_n492_));
  INV_X1    g291(.A(G197gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(G204gat), .ZN(new_n494_));
  INV_X1    g293(.A(G204gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(G204gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n489_), .A2(G211gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n487_), .A2(G218gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n491_), .A2(new_n498_), .A3(KEYINPUT21), .A4(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT21), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n494_), .A2(new_n496_), .A3(new_n504_), .A4(new_n497_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n493_), .A2(G204gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n495_), .A2(G197gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT21), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n488_), .A2(new_n490_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n486_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT29), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n514_), .B2(new_n460_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  OAI221_X1 g315(.A(new_n511_), .B1(new_n512_), .B2(new_n486_), .C1(new_n514_), .C2(new_n460_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n483_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n517_), .A3(new_n483_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n517_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n483_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n482_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT98), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n520_), .A2(new_n519_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n523_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n524_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT98), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n482_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n482_), .A2(new_n518_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n527_), .A2(new_n533_), .B1(new_n520_), .B2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G8gat), .B(G36gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT18), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G64gat), .B(G92gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G226gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT19), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n391_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT22), .B(G169gat), .ZN(new_n545_));
  INV_X1    g344(.A(G176gat), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n410_), .B2(new_n384_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n401_), .A2(new_n403_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n395_), .A2(new_n397_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n392_), .B(new_n383_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT103), .ZN(new_n553_));
  INV_X1    g352(.A(new_n511_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT103), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n555_), .A3(new_n551_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n411_), .B2(new_n511_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n543_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT20), .B1(new_n411_), .B2(new_n511_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n548_), .A2(new_n551_), .B1(new_n510_), .B2(new_n503_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n561_), .A2(new_n542_), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n540_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n542_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n548_), .A2(new_n510_), .A3(new_n503_), .A4(new_n551_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n543_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n539_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(KEYINPUT27), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT27), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n565_), .A2(new_n539_), .A3(new_n567_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n539_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n535_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n474_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n430_), .B(new_n431_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n534_), .A2(new_n520_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n532_), .B1(new_n531_), .B2(new_n482_), .ZN(new_n580_));
  AOI211_X1 g379(.A(KEYINPUT98), .B(new_n481_), .C1(new_n530_), .C2(new_n524_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n539_), .A2(KEYINPUT32), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n565_), .A2(new_n567_), .A3(new_n583_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n585_), .B(new_n586_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT24), .ZN(new_n590_));
  INV_X1    g389(.A(G169gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n546_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n544_), .B2(new_n389_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n399_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n550_), .A2(KEYINPUT88), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n410_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n596_), .A2(new_n597_), .B1(new_n386_), .B2(new_n378_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n558_), .B1(new_n598_), .B2(new_n554_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n562_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n543_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n411_), .A2(new_n511_), .ZN(new_n602_));
  AND4_X1   g401(.A1(KEYINPUT20), .A2(new_n602_), .A3(new_n543_), .A4(new_n566_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n540_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(KEYINPUT99), .A3(new_n568_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n459_), .A2(new_n461_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(KEYINPUT102), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(KEYINPUT102), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n435_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n462_), .A2(new_n435_), .A3(new_n463_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n470_), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n589_), .A2(new_n605_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n472_), .A2(new_n613_), .ZN(new_n614_));
  AOI211_X1 g413(.A(KEYINPUT33), .B(new_n470_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n587_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n578_), .B1(new_n582_), .B2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n569_), .A2(new_n473_), .A3(new_n573_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n527_), .A2(new_n533_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n620_), .B2(new_n579_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT104), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n473_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n582_), .B1(new_n623_), .B2(new_n574_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n472_), .B(new_n613_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n625_), .A2(new_n605_), .A3(new_n611_), .A4(new_n589_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n535_), .A2(new_n587_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n624_), .A2(new_n627_), .A3(new_n628_), .A4(new_n578_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n577_), .B1(new_n622_), .B2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G113gat), .B(G141gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(G169gat), .B(G197gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT87), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n302_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n251_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT85), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n637_), .A2(new_n638_), .B1(new_n302_), .B2(new_n248_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n251_), .A2(KEYINPUT85), .A3(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n639_), .A2(new_n640_), .A3(KEYINPUT86), .A4(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n302_), .B(new_n248_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT84), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(KEYINPUT84), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n637_), .A2(new_n638_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n302_), .A2(new_n248_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n640_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT86), .B1(new_n651_), .B2(new_n641_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n635_), .B1(new_n648_), .B2(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n646_), .A2(new_n647_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n635_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n639_), .A2(new_n641_), .A3(new_n640_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT86), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n654_), .A2(new_n655_), .A3(new_n658_), .A4(new_n642_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n653_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n376_), .A2(new_n630_), .A3(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n329_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(new_n623_), .A3(new_n293_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT105), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n374_), .A2(KEYINPUT13), .A3(new_n368_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT13), .B1(new_n374_), .B2(new_n368_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n660_), .A3(new_n327_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n577_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n587_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n589_), .A2(new_n605_), .A3(new_n611_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n625_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n433_), .B1(new_n675_), .B2(new_n535_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n628_), .B1(new_n676_), .B2(new_n624_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n618_), .A2(KEYINPUT104), .A3(new_n621_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n672_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(KEYINPUT106), .A3(new_n291_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681_));
  INV_X1    g480(.A(new_n291_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n630_), .B2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n671_), .B1(new_n680_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n623_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n664_), .A2(new_n665_), .B1(G1gat), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n667_), .A2(new_n686_), .ZN(G1324gat));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  INV_X1    g487(.A(new_n671_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n680_), .A2(new_n683_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n574_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G8gat), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(KEYINPUT39), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n663_), .A2(new_n294_), .A3(new_n574_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n694_), .B2(KEYINPUT39), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n688_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n694_), .A2(KEYINPUT39), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n701_), .A2(KEYINPUT40), .A3(new_n696_), .A4(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1325gat));
  NAND3_X1  g502(.A1(new_n663_), .A2(new_n417_), .A3(new_n433_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n684_), .A2(new_n433_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT41), .B1(new_n705_), .B2(G15gat), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n707_), .B(new_n417_), .C1(new_n684_), .C2(new_n433_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1326gat));
  INV_X1    g510(.A(G22gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n684_), .B2(new_n582_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT42), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n663_), .A2(new_n712_), .A3(new_n582_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1327gat));
  NOR2_X1   g515(.A1(new_n327_), .A2(new_n291_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n662_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G29gat), .B1(new_n718_), .B2(new_n623_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n279_), .A2(new_n285_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT76), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n279_), .A2(new_n285_), .A3(KEYINPUT76), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n723_), .A2(new_n724_), .B1(new_n682_), .B2(new_n202_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n679_), .A2(new_n720_), .A3(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n630_), .B2(new_n292_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n376_), .A2(new_n661_), .A3(new_n327_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT44), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n623_), .A2(G29gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n719_), .B1(new_n731_), .B2(new_n732_), .ZN(G1328gat));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n575_), .A2(G36gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n718_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT45), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n718_), .A2(new_n739_), .A3(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n731_), .A2(new_n574_), .ZN(new_n741_));
  AOI221_X4 g540(.A(new_n735_), .B1(new_n738_), .B2(new_n740_), .C1(new_n741_), .C2(G36gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(G36gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n738_), .A2(new_n740_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n734_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1329gat));
  AOI21_X1  g545(.A(G43gat), .B1(new_n718_), .B2(new_n433_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT110), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n731_), .A2(G43gat), .A3(new_n433_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT47), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n752_), .A3(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1330gat));
  INV_X1    g553(.A(G50gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n718_), .A2(new_n755_), .A3(new_n582_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n731_), .A2(new_n582_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G50gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT111), .B(new_n755_), .C1(new_n731_), .C2(new_n582_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1331gat));
  INV_X1    g560(.A(G57gat), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n329_), .A2(new_n376_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT112), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n630_), .A2(new_n660_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n329_), .A2(new_n766_), .A3(new_n376_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n768_), .B2(new_n473_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT113), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n762_), .C1(new_n768_), .C2(new_n473_), .ZN(new_n772_));
  AND4_X1   g571(.A1(new_n661_), .A2(new_n690_), .A3(new_n376_), .A4(new_n327_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n473_), .A2(new_n762_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n770_), .A2(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(G1332gat));
  INV_X1    g574(.A(new_n768_), .ZN(new_n776_));
  INV_X1    g575(.A(G64gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n574_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n773_), .A2(new_n574_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G64gat), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT48), .B(new_n777_), .C1(new_n773_), .C2(new_n574_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1333gat));
  INV_X1    g582(.A(G71gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n776_), .A2(new_n784_), .A3(new_n433_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n773_), .A2(new_n433_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(G71gat), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT49), .B(new_n784_), .C1(new_n773_), .C2(new_n433_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1334gat));
  INV_X1    g589(.A(G78gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n776_), .A2(new_n791_), .A3(new_n582_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n773_), .A2(new_n582_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G78gat), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT50), .B(new_n791_), .C1(new_n773_), .C2(new_n582_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(G1335gat));
  AND3_X1   g596(.A1(new_n765_), .A2(new_n376_), .A3(new_n717_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n221_), .A3(new_n623_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n326_), .A2(new_n661_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n727_), .A2(new_n726_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n800_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT114), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT115), .Z(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n623_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n799_), .B1(new_n809_), .B2(new_n221_), .ZN(G1336gat));
  AOI21_X1  g609(.A(G92gat), .B1(new_n798_), .B2(new_n574_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n575_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n808_), .B2(new_n812_), .ZN(G1337gat));
  NAND3_X1  g612(.A1(new_n803_), .A2(new_n433_), .A3(new_n806_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n433_), .A2(new_n236_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n814_), .A2(G99gat), .B1(new_n798_), .B2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n818_), .B(new_n819_), .Z(G1338gat));
  NAND3_X1  g619(.A1(new_n798_), .A2(new_n582_), .A3(new_n237_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n801_), .A2(new_n802_), .ZN(new_n823_));
  AND4_X1   g622(.A1(new_n582_), .A2(new_n728_), .A3(new_n806_), .A4(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n211_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n728_), .A2(new_n806_), .A3(new_n823_), .A4(new_n582_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT117), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n822_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n803_), .A2(new_n825_), .A3(new_n582_), .A4(new_n806_), .ZN(new_n830_));
  AND4_X1   g629(.A1(new_n822_), .A2(new_n828_), .A3(G106gat), .A4(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n821_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT53), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n821_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1339gat));
  NAND2_X1  g635(.A1(new_n370_), .A2(new_n660_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n347_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n354_), .A2(new_n349_), .A3(new_n334_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n840_), .A2(KEYINPUT55), .B1(new_n841_), .B2(new_n336_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n348_), .A2(new_n843_), .A3(new_n356_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n362_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT56), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n370_), .A2(new_n660_), .A3(KEYINPUT118), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n839_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n654_), .A2(new_n633_), .A3(new_n658_), .A4(new_n642_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n651_), .A2(new_n644_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n633_), .B1(new_n643_), .B2(new_n641_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(KEYINPUT119), .A3(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n374_), .B2(new_n368_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n848_), .B1(new_n857_), .B2(KEYINPUT120), .ZN(new_n858_));
  INV_X1    g657(.A(new_n856_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n291_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n845_), .B(KEYINPUT56), .Z(new_n867_));
  NAND2_X1  g666(.A1(new_n859_), .A2(new_n370_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n846_), .A2(KEYINPUT58), .A3(new_n370_), .A4(new_n859_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n725_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n860_), .A2(new_n861_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n857_), .A2(KEYINPUT120), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n848_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n682_), .A2(new_n864_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n871_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n327_), .B1(new_n865_), .B2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n725_), .A2(new_n326_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n670_), .A2(new_n878_), .A3(new_n661_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n877_), .A2(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n576_), .A2(new_n473_), .A3(new_n578_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(G113gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n660_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n871_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n858_), .A2(new_n862_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n875_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n874_), .B2(new_n291_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n326_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n879_), .B(KEYINPUT54), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(KEYINPUT59), .A3(new_n883_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n661_), .B1(new_n889_), .B2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n887_), .B1(new_n899_), .B2(new_n886_), .ZN(G1340gat));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n901_));
  AOI21_X1  g700(.A(G120gat), .B1(new_n376_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT121), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n901_), .B2(G120gat), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n885_), .B(new_n903_), .C1(new_n902_), .C2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n670_), .B1(new_n889_), .B2(new_n898_), .ZN(new_n907_));
  INV_X1    g706(.A(G120gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1341gat));
  OAI211_X1 g708(.A(new_n327_), .B(new_n883_), .C1(new_n877_), .C2(new_n881_), .ZN(new_n910_));
  INV_X1    g709(.A(G127gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT122), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n910_), .A2(new_n914_), .A3(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n889_), .A2(new_n898_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n326_), .A2(new_n911_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n913_), .A2(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1342gat));
  INV_X1    g717(.A(G134gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n885_), .A2(new_n919_), .A3(new_n682_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n292_), .B1(new_n889_), .B2(new_n898_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n919_), .ZN(G1343gat));
  NOR4_X1   g721(.A1(new_n433_), .A2(new_n535_), .A3(new_n473_), .A4(new_n574_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n897_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n660_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(G141gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n438_), .A3(new_n660_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1344gat));
  NAND2_X1  g727(.A1(new_n924_), .A2(new_n376_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G148gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n924_), .A2(new_n439_), .A3(new_n376_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1345gat));
  OAI211_X1 g731(.A(new_n327_), .B(new_n923_), .C1(new_n877_), .C2(new_n881_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(KEYINPUT123), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n897_), .A2(new_n935_), .A3(new_n327_), .A4(new_n923_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT61), .B(G155gat), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n934_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1346gat));
  NAND2_X1  g739(.A1(new_n924_), .A2(new_n682_), .ZN(new_n941_));
  INV_X1    g740(.A(G162gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n725_), .A2(G162gat), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n943_), .B(KEYINPUT124), .Z(new_n944_));
  AOI22_X1  g743(.A1(new_n941_), .A2(new_n942_), .B1(new_n924_), .B2(new_n944_), .ZN(G1347gat));
  NOR3_X1   g744(.A1(new_n474_), .A2(new_n582_), .A3(new_n575_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n897_), .A2(new_n660_), .A3(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(G169gat), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n897_), .A2(new_n946_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n951_), .A2(new_n545_), .A3(new_n660_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n947_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n950_), .A2(new_n952_), .A3(new_n953_), .ZN(G1348gat));
  NAND3_X1  g753(.A1(new_n897_), .A2(new_n376_), .A3(new_n946_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g755(.A1(new_n897_), .A2(new_n327_), .A3(new_n946_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n550_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n959_), .B1(new_n396_), .B2(new_n957_), .ZN(G1350gat));
  NAND4_X1  g759(.A1(new_n951_), .A2(new_n401_), .A3(new_n403_), .A4(new_n682_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n897_), .A2(new_n725_), .A3(new_n946_), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n962_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n963_));
  AOI21_X1  g762(.A(KEYINPUT125), .B1(new_n962_), .B2(G190gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n961_), .B1(new_n963_), .B2(new_n964_), .ZN(G1351gat));
  NOR4_X1   g764(.A1(new_n433_), .A2(new_n535_), .A3(new_n623_), .A4(new_n575_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n660_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n376_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(KEYINPUT126), .ZN(new_n974_));
  NAND2_X1  g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  NAND4_X1  g774(.A1(new_n968_), .A2(new_n327_), .A3(new_n974_), .A4(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n973_), .A2(KEYINPUT126), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n976_), .B(new_n977_), .ZN(G1354gat));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n489_), .B1(new_n968_), .B2(new_n725_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n682_), .A2(new_n489_), .ZN(new_n981_));
  NOR3_X1   g780(.A1(new_n882_), .A2(new_n967_), .A3(new_n981_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n979_), .B1(new_n980_), .B2(new_n982_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n968_), .A2(new_n489_), .A3(new_n682_), .ZN(new_n984_));
  NOR3_X1   g783(.A1(new_n882_), .A2(new_n292_), .A3(new_n967_), .ZN(new_n985_));
  OAI211_X1 g784(.A(KEYINPUT127), .B(new_n984_), .C1(new_n985_), .C2(new_n489_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n983_), .A2(new_n986_), .ZN(G1355gat));
endmodule


